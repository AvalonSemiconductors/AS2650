magic
tech gf180mcuC
magscale 1 5
timestamp 1670429284
<< obsm1 >>
rect 672 1538 89320 58561
<< metal2 >>
rect 672 59600 728 60000
rect 1456 59600 1512 60000
rect 2240 59600 2296 60000
rect 3024 59600 3080 60000
rect 3808 59600 3864 60000
rect 4592 59600 4648 60000
rect 5376 59600 5432 60000
rect 6160 59600 6216 60000
rect 6944 59600 7000 60000
rect 7728 59600 7784 60000
rect 8512 59600 8568 60000
rect 9296 59600 9352 60000
rect 10080 59600 10136 60000
rect 10864 59600 10920 60000
rect 11648 59600 11704 60000
rect 12432 59600 12488 60000
rect 13216 59600 13272 60000
rect 14000 59600 14056 60000
rect 14784 59600 14840 60000
rect 15568 59600 15624 60000
rect 16352 59600 16408 60000
rect 17136 59600 17192 60000
rect 17920 59600 17976 60000
rect 18704 59600 18760 60000
rect 19488 59600 19544 60000
rect 20272 59600 20328 60000
rect 21056 59600 21112 60000
rect 21840 59600 21896 60000
rect 22624 59600 22680 60000
rect 23408 59600 23464 60000
rect 24192 59600 24248 60000
rect 24976 59600 25032 60000
rect 25760 59600 25816 60000
rect 26544 59600 26600 60000
rect 27328 59600 27384 60000
rect 28112 59600 28168 60000
rect 28896 59600 28952 60000
rect 29680 59600 29736 60000
rect 30464 59600 30520 60000
rect 31248 59600 31304 60000
rect 32032 59600 32088 60000
rect 32816 59600 32872 60000
rect 33600 59600 33656 60000
rect 34384 59600 34440 60000
rect 35168 59600 35224 60000
rect 35952 59600 36008 60000
rect 36736 59600 36792 60000
rect 37520 59600 37576 60000
rect 38304 59600 38360 60000
rect 39088 59600 39144 60000
rect 39872 59600 39928 60000
rect 40656 59600 40712 60000
rect 41440 59600 41496 60000
rect 42224 59600 42280 60000
rect 43008 59600 43064 60000
rect 43792 59600 43848 60000
rect 44576 59600 44632 60000
rect 45360 59600 45416 60000
rect 46144 59600 46200 60000
rect 46928 59600 46984 60000
rect 47712 59600 47768 60000
rect 48496 59600 48552 60000
rect 49280 59600 49336 60000
rect 50064 59600 50120 60000
rect 50848 59600 50904 60000
rect 51632 59600 51688 60000
rect 52416 59600 52472 60000
rect 53200 59600 53256 60000
rect 53984 59600 54040 60000
rect 54768 59600 54824 60000
rect 55552 59600 55608 60000
rect 56336 59600 56392 60000
rect 57120 59600 57176 60000
rect 57904 59600 57960 60000
rect 58688 59600 58744 60000
rect 59472 59600 59528 60000
rect 60256 59600 60312 60000
rect 61040 59600 61096 60000
rect 61824 59600 61880 60000
rect 62608 59600 62664 60000
rect 63392 59600 63448 60000
rect 64176 59600 64232 60000
rect 64960 59600 65016 60000
rect 65744 59600 65800 60000
rect 66528 59600 66584 60000
rect 67312 59600 67368 60000
rect 68096 59600 68152 60000
rect 68880 59600 68936 60000
rect 69664 59600 69720 60000
rect 70448 59600 70504 60000
rect 71232 59600 71288 60000
rect 72016 59600 72072 60000
rect 72800 59600 72856 60000
rect 73584 59600 73640 60000
rect 74368 59600 74424 60000
rect 75152 59600 75208 60000
rect 75936 59600 75992 60000
rect 76720 59600 76776 60000
rect 77504 59600 77560 60000
rect 78288 59600 78344 60000
rect 79072 59600 79128 60000
rect 79856 59600 79912 60000
rect 80640 59600 80696 60000
rect 81424 59600 81480 60000
rect 82208 59600 82264 60000
rect 82992 59600 83048 60000
rect 83776 59600 83832 60000
rect 84560 59600 84616 60000
rect 85344 59600 85400 60000
rect 86128 59600 86184 60000
rect 86912 59600 86968 60000
rect 87696 59600 87752 60000
rect 88480 59600 88536 60000
rect 89264 59600 89320 60000
rect 22456 0 22512 400
rect 67424 0 67480 400
<< obsm2 >>
rect 758 59570 1426 59855
rect 1542 59570 2210 59855
rect 2326 59570 2994 59855
rect 3110 59570 3778 59855
rect 3894 59570 4562 59855
rect 4678 59570 5346 59855
rect 5462 59570 6130 59855
rect 6246 59570 6914 59855
rect 7030 59570 7698 59855
rect 7814 59570 8482 59855
rect 8598 59570 9266 59855
rect 9382 59570 10050 59855
rect 10166 59570 10834 59855
rect 10950 59570 11618 59855
rect 11734 59570 12402 59855
rect 12518 59570 13186 59855
rect 13302 59570 13970 59855
rect 14086 59570 14754 59855
rect 14870 59570 15538 59855
rect 15654 59570 16322 59855
rect 16438 59570 17106 59855
rect 17222 59570 17890 59855
rect 18006 59570 18674 59855
rect 18790 59570 19458 59855
rect 19574 59570 20242 59855
rect 20358 59570 21026 59855
rect 21142 59570 21810 59855
rect 21926 59570 22594 59855
rect 22710 59570 23378 59855
rect 23494 59570 24162 59855
rect 24278 59570 24946 59855
rect 25062 59570 25730 59855
rect 25846 59570 26514 59855
rect 26630 59570 27298 59855
rect 27414 59570 28082 59855
rect 28198 59570 28866 59855
rect 28982 59570 29650 59855
rect 29766 59570 30434 59855
rect 30550 59570 31218 59855
rect 31334 59570 32002 59855
rect 32118 59570 32786 59855
rect 32902 59570 33570 59855
rect 33686 59570 34354 59855
rect 34470 59570 35138 59855
rect 35254 59570 35922 59855
rect 36038 59570 36706 59855
rect 36822 59570 37490 59855
rect 37606 59570 38274 59855
rect 38390 59570 39058 59855
rect 39174 59570 39842 59855
rect 39958 59570 40626 59855
rect 40742 59570 41410 59855
rect 41526 59570 42194 59855
rect 42310 59570 42978 59855
rect 43094 59570 43762 59855
rect 43878 59570 44546 59855
rect 44662 59570 45330 59855
rect 45446 59570 46114 59855
rect 46230 59570 46898 59855
rect 47014 59570 47682 59855
rect 47798 59570 48466 59855
rect 48582 59570 49250 59855
rect 49366 59570 50034 59855
rect 50150 59570 50818 59855
rect 50934 59570 51602 59855
rect 51718 59570 52386 59855
rect 52502 59570 53170 59855
rect 53286 59570 53954 59855
rect 54070 59570 54738 59855
rect 54854 59570 55522 59855
rect 55638 59570 56306 59855
rect 56422 59570 57090 59855
rect 57206 59570 57874 59855
rect 57990 59570 58658 59855
rect 58774 59570 59442 59855
rect 59558 59570 60226 59855
rect 60342 59570 61010 59855
rect 61126 59570 61794 59855
rect 61910 59570 62578 59855
rect 62694 59570 63362 59855
rect 63478 59570 64146 59855
rect 64262 59570 64930 59855
rect 65046 59570 65714 59855
rect 65830 59570 66498 59855
rect 66614 59570 67282 59855
rect 67398 59570 68066 59855
rect 68182 59570 68850 59855
rect 68966 59570 69634 59855
rect 69750 59570 70418 59855
rect 70534 59570 71202 59855
rect 71318 59570 71986 59855
rect 72102 59570 72770 59855
rect 72886 59570 73554 59855
rect 73670 59570 74338 59855
rect 74454 59570 75122 59855
rect 75238 59570 75906 59855
rect 76022 59570 76690 59855
rect 76806 59570 77474 59855
rect 77590 59570 78258 59855
rect 78374 59570 79042 59855
rect 79158 59570 79826 59855
rect 79942 59570 80610 59855
rect 80726 59570 81394 59855
rect 81510 59570 82178 59855
rect 82294 59570 82962 59855
rect 83078 59570 83746 59855
rect 83862 59570 84530 59855
rect 84646 59570 85314 59855
rect 85430 59570 86098 59855
rect 86214 59570 86882 59855
rect 86998 59570 87666 59855
rect 87782 59570 88450 59855
rect 88566 59570 89234 59855
rect 742 430 89306 59570
rect 742 400 22426 430
rect 22542 400 67394 430
rect 67510 400 89306 430
<< obsm3 >>
rect 737 1302 89311 59850
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
rect 86704 1538 86864 58438
<< obsm4 >>
rect 4158 58468 86954 59015
rect 4158 1508 9874 58468
rect 10094 1508 17554 58468
rect 17774 1508 25234 58468
rect 25454 1508 32914 58468
rect 33134 1508 40594 58468
rect 40814 1508 48274 58468
rect 48494 1508 55954 58468
rect 56174 1508 63634 58468
rect 63854 1508 71314 58468
rect 71534 1508 78994 58468
rect 79214 1508 86674 58468
rect 86894 1508 86954 58468
rect 4158 1297 86954 1508
<< labels >>
rlabel metal2 s 672 59600 728 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24192 59600 24248 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 26544 59600 26600 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 28896 59600 28952 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 31248 59600 31304 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 33600 59600 33656 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 35952 59600 36008 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 38304 59600 38360 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 40656 59600 40712 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 43008 59600 43064 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 45360 59600 45416 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3024 59600 3080 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 47712 59600 47768 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 50064 59600 50120 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 52416 59600 52472 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 54768 59600 54824 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 57120 59600 57176 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 59472 59600 59528 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 61824 59600 61880 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 64176 59600 64232 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 66528 59600 66584 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 68880 59600 68936 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5376 59600 5432 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 71232 59600 71288 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 73584 59600 73640 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 75936 59600 75992 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 78288 59600 78344 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 80640 59600 80696 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 82992 59600 83048 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 85344 59600 85400 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 87696 59600 87752 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7728 59600 7784 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10080 59600 10136 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 12432 59600 12488 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 14784 59600 14840 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 17136 59600 17192 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 19488 59600 19544 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 21840 59600 21896 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1456 59600 1512 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 24976 59600 25032 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 27328 59600 27384 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 29680 59600 29736 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 32032 59600 32088 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 34384 59600 34440 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 36736 59600 36792 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 39088 59600 39144 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 41440 59600 41496 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 43792 59600 43848 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 46144 59600 46200 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3808 59600 3864 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 48496 59600 48552 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 50848 59600 50904 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 53200 59600 53256 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 55552 59600 55608 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 57904 59600 57960 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 60256 59600 60312 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 62608 59600 62664 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 64960 59600 65016 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 67312 59600 67368 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 69664 59600 69720 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6160 59600 6216 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 72016 59600 72072 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 74368 59600 74424 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 76720 59600 76776 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 79072 59600 79128 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 81424 59600 81480 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 83776 59600 83832 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 86128 59600 86184 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 88480 59600 88536 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8512 59600 8568 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10864 59600 10920 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13216 59600 13272 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 15568 59600 15624 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 17920 59600 17976 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 20272 59600 20328 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 22624 59600 22680 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2240 59600 2296 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 25760 59600 25816 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 28112 59600 28168 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 30464 59600 30520 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 32816 59600 32872 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 35168 59600 35224 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 37520 59600 37576 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 39872 59600 39928 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 42224 59600 42280 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 44576 59600 44632 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 46928 59600 46984 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4592 59600 4648 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 49280 59600 49336 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 51632 59600 51688 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 53984 59600 54040 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 56336 59600 56392 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 58688 59600 58744 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 61040 59600 61096 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 63392 59600 63448 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 65744 59600 65800 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 68096 59600 68152 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 70448 59600 70504 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 6944 59600 7000 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 72800 59600 72856 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 75152 59600 75208 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 77504 59600 77560 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 79856 59600 79912 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 82208 59600 82264 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 84560 59600 84616 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 86912 59600 86968 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 89264 59600 89320 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9296 59600 9352 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11648 59600 11704 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14000 59600 14056 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 16352 59600 16408 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 18704 59600 18760 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 21056 59600 21112 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 23408 59600 23464 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 58438 6 vss
port 116 nsew ground bidirectional
rlabel metal2 s 22456 0 22512 400 6 wb_clk_i
port 117 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 wb_rst_i
port 118 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12724232
string GDS_FILE /home/lucah/Videos/AS2650/openlane/wrapped_as2650/runs/22_12_07_17_02/results/signoff/wrapped_as2650.magic.gds
string GDS_START 387682
<< end >>

