// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 output [63:0] la_data_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire net194;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net197;
 wire net145;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net146;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net195;
 wire net196;
 wire net153;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net154;
 wire net155;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire \as2650.PC[0] ;
 wire \as2650.PC[10] ;
 wire \as2650.PC[11] ;
 wire \as2650.PC[12] ;
 wire \as2650.PC[1] ;
 wire \as2650.PC[2] ;
 wire \as2650.PC[3] ;
 wire \as2650.PC[4] ;
 wire \as2650.PC[5] ;
 wire \as2650.PC[6] ;
 wire \as2650.PC[7] ;
 wire \as2650.PC[8] ;
 wire \as2650.PC[9] ;
 wire \as2650.chirp_ptr[0] ;
 wire \as2650.chirp_ptr[1] ;
 wire \as2650.chirp_ptr[2] ;
 wire \as2650.chirpchar[0] ;
 wire \as2650.chirpchar[1] ;
 wire \as2650.chirpchar[2] ;
 wire \as2650.chirpchar[3] ;
 wire \as2650.chirpchar[4] ;
 wire \as2650.chirpchar[5] ;
 wire \as2650.chirpchar[6] ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.debug_psl[0] ;
 wire \as2650.debug_psl[1] ;
 wire \as2650.debug_psl[2] ;
 wire \as2650.debug_psl[3] ;
 wire \as2650.debug_psl[4] ;
 wire \as2650.debug_psl[5] ;
 wire \as2650.debug_psl[6] ;
 wire \as2650.debug_psl[7] ;
 wire \as2650.debug_psu[0] ;
 wire \as2650.debug_psu[1] ;
 wire \as2650.debug_psu[2] ;
 wire \as2650.debug_psu[3] ;
 wire \as2650.debug_psu[4] ;
 wire \as2650.debug_psu[5] ;
 wire \as2650.debug_psu[7] ;
 wire \as2650.extend ;
 wire \as2650.indexed_cyc[0] ;
 wire \as2650.indexed_cyc[1] ;
 wire \as2650.indirect_cyc ;
 wire \as2650.indirect_target[0] ;
 wire \as2650.indirect_target[10] ;
 wire \as2650.indirect_target[11] ;
 wire \as2650.indirect_target[12] ;
 wire \as2650.indirect_target[13] ;
 wire \as2650.indirect_target[14] ;
 wire \as2650.indirect_target[15] ;
 wire \as2650.indirect_target[1] ;
 wire \as2650.indirect_target[2] ;
 wire \as2650.indirect_target[3] ;
 wire \as2650.indirect_target[4] ;
 wire \as2650.indirect_target[5] ;
 wire \as2650.indirect_target[6] ;
 wire \as2650.indirect_target[7] ;
 wire \as2650.indirect_target[8] ;
 wire \as2650.indirect_target[9] ;
 wire \as2650.insin[0] ;
 wire \as2650.insin[1] ;
 wire \as2650.insin[2] ;
 wire \as2650.insin[3] ;
 wire \as2650.insin[4] ;
 wire \as2650.insin[5] ;
 wire \as2650.insin[6] ;
 wire \as2650.insin[7] ;
 wire \as2650.instruction_args_latch[0] ;
 wire \as2650.instruction_args_latch[10] ;
 wire \as2650.instruction_args_latch[11] ;
 wire \as2650.instruction_args_latch[12] ;
 wire \as2650.instruction_args_latch[13] ;
 wire \as2650.instruction_args_latch[14] ;
 wire \as2650.instruction_args_latch[15] ;
 wire \as2650.instruction_args_latch[1] ;
 wire \as2650.instruction_args_latch[2] ;
 wire \as2650.instruction_args_latch[3] ;
 wire \as2650.instruction_args_latch[4] ;
 wire \as2650.instruction_args_latch[5] ;
 wire \as2650.instruction_args_latch[6] ;
 wire \as2650.instruction_args_latch[7] ;
 wire \as2650.instruction_args_latch[8] ;
 wire \as2650.instruction_args_latch[9] ;
 wire \as2650.last_addr[0] ;
 wire \as2650.last_addr[10] ;
 wire \as2650.last_addr[11] ;
 wire \as2650.last_addr[12] ;
 wire \as2650.last_addr[13] ;
 wire \as2650.last_addr[14] ;
 wire \as2650.last_addr[15] ;
 wire \as2650.last_addr[1] ;
 wire \as2650.last_addr[2] ;
 wire \as2650.last_addr[3] ;
 wire \as2650.last_addr[4] ;
 wire \as2650.last_addr[5] ;
 wire \as2650.last_addr[6] ;
 wire \as2650.last_addr[7] ;
 wire \as2650.last_addr[8] ;
 wire \as2650.last_addr[9] ;
 wire \as2650.page_reg[0] ;
 wire \as2650.page_reg[1] ;
 wire \as2650.page_reg[2] ;
 wire \as2650.regs[0][0] ;
 wire \as2650.regs[0][1] ;
 wire \as2650.regs[0][2] ;
 wire \as2650.regs[0][3] ;
 wire \as2650.regs[0][4] ;
 wire \as2650.regs[0][5] ;
 wire \as2650.regs[0][6] ;
 wire \as2650.regs[0][7] ;
 wire \as2650.regs[1][0] ;
 wire \as2650.regs[1][1] ;
 wire \as2650.regs[1][2] ;
 wire \as2650.regs[1][3] ;
 wire \as2650.regs[1][4] ;
 wire \as2650.regs[1][5] ;
 wire \as2650.regs[1][6] ;
 wire \as2650.regs[1][7] ;
 wire \as2650.regs[2][0] ;
 wire \as2650.regs[2][1] ;
 wire \as2650.regs[2][2] ;
 wire \as2650.regs[2][3] ;
 wire \as2650.regs[2][4] ;
 wire \as2650.regs[2][5] ;
 wire \as2650.regs[2][6] ;
 wire \as2650.regs[2][7] ;
 wire \as2650.regs[3][0] ;
 wire \as2650.regs[3][1] ;
 wire \as2650.regs[3][2] ;
 wire \as2650.regs[3][3] ;
 wire \as2650.regs[3][4] ;
 wire \as2650.regs[3][5] ;
 wire \as2650.regs[3][6] ;
 wire \as2650.regs[3][7] ;
 wire \as2650.regs[4][0] ;
 wire \as2650.regs[4][1] ;
 wire \as2650.regs[4][2] ;
 wire \as2650.regs[4][3] ;
 wire \as2650.regs[4][4] ;
 wire \as2650.regs[4][5] ;
 wire \as2650.regs[4][6] ;
 wire \as2650.regs[4][7] ;
 wire \as2650.regs[5][0] ;
 wire \as2650.regs[5][1] ;
 wire \as2650.regs[5][2] ;
 wire \as2650.regs[5][3] ;
 wire \as2650.regs[5][4] ;
 wire \as2650.regs[5][5] ;
 wire \as2650.regs[5][6] ;
 wire \as2650.regs[5][7] ;
 wire \as2650.regs[6][0] ;
 wire \as2650.regs[6][1] ;
 wire \as2650.regs[6][2] ;
 wire \as2650.regs[6][3] ;
 wire \as2650.regs[6][4] ;
 wire \as2650.regs[6][5] ;
 wire \as2650.regs[6][6] ;
 wire \as2650.regs[6][7] ;
 wire \as2650.regs[7][0] ;
 wire \as2650.regs[7][1] ;
 wire \as2650.regs[7][2] ;
 wire \as2650.regs[7][3] ;
 wire \as2650.regs[7][4] ;
 wire \as2650.regs[7][5] ;
 wire \as2650.regs[7][6] ;
 wire \as2650.regs[7][7] ;
 wire \as2650.relative_cyc ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][15] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[10][0] ;
 wire \as2650.stack[10][10] ;
 wire \as2650.stack[10][11] ;
 wire \as2650.stack[10][12] ;
 wire \as2650.stack[10][13] ;
 wire \as2650.stack[10][14] ;
 wire \as2650.stack[10][15] ;
 wire \as2650.stack[10][1] ;
 wire \as2650.stack[10][2] ;
 wire \as2650.stack[10][3] ;
 wire \as2650.stack[10][4] ;
 wire \as2650.stack[10][5] ;
 wire \as2650.stack[10][6] ;
 wire \as2650.stack[10][7] ;
 wire \as2650.stack[10][8] ;
 wire \as2650.stack[10][9] ;
 wire \as2650.stack[11][0] ;
 wire \as2650.stack[11][10] ;
 wire \as2650.stack[11][11] ;
 wire \as2650.stack[11][12] ;
 wire \as2650.stack[11][13] ;
 wire \as2650.stack[11][14] ;
 wire \as2650.stack[11][15] ;
 wire \as2650.stack[11][1] ;
 wire \as2650.stack[11][2] ;
 wire \as2650.stack[11][3] ;
 wire \as2650.stack[11][4] ;
 wire \as2650.stack[11][5] ;
 wire \as2650.stack[11][6] ;
 wire \as2650.stack[11][7] ;
 wire \as2650.stack[11][8] ;
 wire \as2650.stack[11][9] ;
 wire \as2650.stack[12][0] ;
 wire \as2650.stack[12][10] ;
 wire \as2650.stack[12][11] ;
 wire \as2650.stack[12][12] ;
 wire \as2650.stack[12][13] ;
 wire \as2650.stack[12][14] ;
 wire \as2650.stack[12][15] ;
 wire \as2650.stack[12][1] ;
 wire \as2650.stack[12][2] ;
 wire \as2650.stack[12][3] ;
 wire \as2650.stack[12][4] ;
 wire \as2650.stack[12][5] ;
 wire \as2650.stack[12][6] ;
 wire \as2650.stack[12][7] ;
 wire \as2650.stack[12][8] ;
 wire \as2650.stack[12][9] ;
 wire \as2650.stack[13][0] ;
 wire \as2650.stack[13][10] ;
 wire \as2650.stack[13][11] ;
 wire \as2650.stack[13][12] ;
 wire \as2650.stack[13][13] ;
 wire \as2650.stack[13][14] ;
 wire \as2650.stack[13][15] ;
 wire \as2650.stack[13][1] ;
 wire \as2650.stack[13][2] ;
 wire \as2650.stack[13][3] ;
 wire \as2650.stack[13][4] ;
 wire \as2650.stack[13][5] ;
 wire \as2650.stack[13][6] ;
 wire \as2650.stack[13][7] ;
 wire \as2650.stack[13][8] ;
 wire \as2650.stack[13][9] ;
 wire \as2650.stack[14][0] ;
 wire \as2650.stack[14][10] ;
 wire \as2650.stack[14][11] ;
 wire \as2650.stack[14][12] ;
 wire \as2650.stack[14][13] ;
 wire \as2650.stack[14][14] ;
 wire \as2650.stack[14][15] ;
 wire \as2650.stack[14][1] ;
 wire \as2650.stack[14][2] ;
 wire \as2650.stack[14][3] ;
 wire \as2650.stack[14][4] ;
 wire \as2650.stack[14][5] ;
 wire \as2650.stack[14][6] ;
 wire \as2650.stack[14][7] ;
 wire \as2650.stack[14][8] ;
 wire \as2650.stack[14][9] ;
 wire \as2650.stack[15][0] ;
 wire \as2650.stack[15][10] ;
 wire \as2650.stack[15][11] ;
 wire \as2650.stack[15][12] ;
 wire \as2650.stack[15][13] ;
 wire \as2650.stack[15][14] ;
 wire \as2650.stack[15][15] ;
 wire \as2650.stack[15][1] ;
 wire \as2650.stack[15][2] ;
 wire \as2650.stack[15][3] ;
 wire \as2650.stack[15][4] ;
 wire \as2650.stack[15][5] ;
 wire \as2650.stack[15][6] ;
 wire \as2650.stack[15][7] ;
 wire \as2650.stack[15][8] ;
 wire \as2650.stack[15][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][15] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][15] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][15] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][15] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][15] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][15] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][15] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack[8][0] ;
 wire \as2650.stack[8][10] ;
 wire \as2650.stack[8][11] ;
 wire \as2650.stack[8][12] ;
 wire \as2650.stack[8][13] ;
 wire \as2650.stack[8][14] ;
 wire \as2650.stack[8][15] ;
 wire \as2650.stack[8][1] ;
 wire \as2650.stack[8][2] ;
 wire \as2650.stack[8][3] ;
 wire \as2650.stack[8][4] ;
 wire \as2650.stack[8][5] ;
 wire \as2650.stack[8][6] ;
 wire \as2650.stack[8][7] ;
 wire \as2650.stack[8][8] ;
 wire \as2650.stack[8][9] ;
 wire \as2650.stack[9][0] ;
 wire \as2650.stack[9][10] ;
 wire \as2650.stack[9][11] ;
 wire \as2650.stack[9][12] ;
 wire \as2650.stack[9][13] ;
 wire \as2650.stack[9][14] ;
 wire \as2650.stack[9][15] ;
 wire \as2650.stack[9][1] ;
 wire \as2650.stack[9][2] ;
 wire \as2650.stack[9][3] ;
 wire \as2650.stack[9][4] ;
 wire \as2650.stack[9][5] ;
 wire \as2650.stack[9][6] ;
 wire \as2650.stack[9][7] ;
 wire \as2650.stack[9][8] ;
 wire \as2650.stack[9][9] ;
 wire \as2650.warmup[0] ;
 wire \as2650.warmup[1] ;
 wire clknet_0__01311_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf__01311_;
 wire clknet_1_1__leaf__01311_;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \wb_counter[0] ;
 wire \wb_counter[10] ;
 wire \wb_counter[11] ;
 wire \wb_counter[12] ;
 wire \wb_counter[13] ;
 wire \wb_counter[14] ;
 wire \wb_counter[15] ;
 wire \wb_counter[16] ;
 wire \wb_counter[17] ;
 wire \wb_counter[18] ;
 wire \wb_counter[19] ;
 wire \wb_counter[1] ;
 wire \wb_counter[20] ;
 wire \wb_counter[21] ;
 wire \wb_counter[22] ;
 wire \wb_counter[23] ;
 wire \wb_counter[24] ;
 wire \wb_counter[25] ;
 wire \wb_counter[26] ;
 wire \wb_counter[27] ;
 wire \wb_counter[28] ;
 wire \wb_counter[29] ;
 wire \wb_counter[2] ;
 wire \wb_counter[30] ;
 wire \wb_counter[31] ;
 wire \wb_counter[3] ;
 wire \wb_counter[4] ;
 wire \wb_counter[5] ;
 wire \wb_counter[6] ;
 wire \wb_counter[7] ;
 wire \wb_counter[8] ;
 wire \wb_counter[9] ;
 wire wb_debug_carry;
 wire wb_debug_cc;
 wire wb_feedback_delay;
 wire \web_behavior[0] ;
 wire \web_behavior[1] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05231__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05232__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05234__I (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05235__I (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05236__I (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05237__I (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05238__I (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05240__I (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05244__I (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05247__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05248__A1 (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05250__I (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05253__I (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05256__A2 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__I (.I(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05258__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05261__I (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05263__I (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05266__A1 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05266__A2 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05267__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05267__A2 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05268__A1 (.I(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05268__A2 (.I(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05269__A1 (.I(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05273__I (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__A2 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__A1 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05280__A2 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05280__B1 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05280__B2 (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05287__B1 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05287__B2 (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05290__B1 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05290__B2 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05293__A1 (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05295__I (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05296__A3 (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05299__A1 (.I(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05299__A2 (.I(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05302__A1 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05302__A2 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05303__A1 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05303__A3 (.I(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05306__A1 (.I(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05307__A2 (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05308__A1 (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05308__A2 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__A2 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__B1 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05310__A1 (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05310__A2 (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__I (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05312__A2 (.I(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05312__B1 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05314__A1 (.I(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05315__I (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__A2 (.I(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05317__A2 (.I(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05319__I (.I(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05324__B2 (.I(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05327__I (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05329__B (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05330__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05331__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05334__A1 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05334__A2 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05336__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05337__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05340__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05343__A1 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05344__B (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__A2 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__B1 (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__B2 (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05348__A1 (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05348__A2 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05352__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05352__A2 (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05352__A3 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__A1 (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05356__A2 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__A2 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05360__A1 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05361__I (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05365__I (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05367__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05368__I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05369__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05371__A1 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05371__A2 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05372__I (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05374__I (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05375__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05377__I (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05380__A2 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05380__B (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05381__A2 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05382__I (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05385__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05386__A2 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05387__I (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05389__I (.I(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05391__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05392__A2 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05393__I (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__B1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__B2 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__C2 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__A1 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__A2 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05402__A2 (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05402__B (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__A1 (.I(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__A2 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__B2 (.I(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05405__A1 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05407__A1 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05408__I (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05410__I (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05411__I (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__A1 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05414__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05415__B (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05416__I (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05417__A1 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05419__A1 (.I(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__A1 (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__A2 (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05422__A1 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__A2 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__B1 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05425__A1 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05426__B (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05427__A1 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05429__A2 (.I(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05431__A1 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05433__C2 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05435__B (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__A1 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__C2 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05438__A1 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05439__I (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05440__B (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05441__B1 (.I(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05441__C2 (.I(\as2650.regs[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05443__B (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__A1 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__B1 (.I(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__C2 (.I(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__A1 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__A2 (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__A1 (.I(\as2650.regs[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__B (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05451__I (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05453__I (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05454__C1 (.I(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05457__A1 (.I(\as2650.regs[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05457__B (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05458__A1 (.I(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05458__C1 (.I(\as2650.regs[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05462__A1 (.I(\as2650.regs[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05462__B (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05463__B1 (.I(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05463__C1 (.I(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05465__I (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05466__A1 (.I(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__A1 (.I(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__C1 (.I(\as2650.regs[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__A1 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__A2 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05472__A1 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05473__C1 (.I(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05473__C2 (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05476__A1 (.I(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05476__B (.I(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__B1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__C1 (.I(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__C2 (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05479__A1 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05481__A1 (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05483__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05483__A2 (.I(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05485__A1 (.I(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__A1 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__A2 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05488__A1 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05488__A2 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__A1 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__A2 (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05490__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05493__A1 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05493__A2 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05495__A1 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__A1 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05501__I (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__A1 (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__A2 (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__B1 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__B2 (.I(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__C1 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__C2 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05507__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05510__A2 (.I(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05513__I (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__A1 (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__A2 (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__A1 (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__A2 (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05520__A3 (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05523__I (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05525__A2 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05526__A1 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05527__I (.I(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05529__A2 (.I(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05530__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05538__A1 (.I(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05541__A2 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__C (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05543__A1 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05544__A1 (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05545__A2 (.I(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__A1 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__A2 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05550__A1 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05552__A1 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05553__A1 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05556__A2 (.I(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05558__B1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05558__B2 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05558__C2 (.I(\as2650.PC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__A1 (.I(\as2650.instruction_args_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05561__A1 (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05561__A2 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05561__A3 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__A1 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__A2 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__A3 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__B (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05565__A2 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05565__B2 (.I(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__A2 (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__B (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05570__A2 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05570__A3 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05574__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05577__A2 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05578__B (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__A1 (.I(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__A2 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__B1 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05582__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05583__A2 (.I(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__A2 (.I(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__A2 (.I(\as2650.instruction_args_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__B (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05588__A4 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05594__A1 (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05595__A1 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05596__A2 (.I(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__A2 (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05601__A2 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05601__A3 (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__A1 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__A1 (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__A2 (.I(\as2650.instruction_args_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__B (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05617__A4 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05618__A2 (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05620__A1 (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05620__A2 (.I(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05623__A2 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05627__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__A2 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__A3 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__B (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__A2 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__A3 (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__B2 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__A2 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__B (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05638__A4 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05639__A2 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05639__A4 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05645__B (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05647__B (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05648__I (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05650__A2 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05652__A1 (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05652__A2 (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05655__A2 (.I(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05656__A1 (.I(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05658__A2 (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__A2 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__A3 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05663__A1 (.I(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__A1 (.I(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__A2 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05665__A1 (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__A2 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05667__I (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05668__A1 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05668__A2 (.I(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05668__B (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05669__B2 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05671__I (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__B1 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__B2 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__A3 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05674__I (.I(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__A1 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__A2 (.I(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05680__A1 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05680__A2 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05682__A1 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05683__A1 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05683__A2 (.I(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05686__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05687__A2 (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05688__A2 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05695__I (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05696__A1 (.I(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__A1 (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05700__A1 (.I(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05704__A1 (.I(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05705__A2 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05707__A1 (.I(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05707__A2 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__A2 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05719__A2 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__A2 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05721__A2 (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05722__A2 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05723__A2 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__A2 (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05725__A2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05726__A2 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05727__A2 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05729__A2 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05730__A2 (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__A2 (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__A2 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05737__A2 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05741__A2 (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__A2 (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__A3 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__A2 (.I(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__I0 (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__I1 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__I (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05749__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__A1 (.I(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__B (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05755__I (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__A1 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__A2 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__B (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__A2 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__A1 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__A2 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__I (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A1 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A2 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__I (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__I (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__A2 (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__I (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__B (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__I (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__A1 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__I (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05776__A1 (.I(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__A2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__I (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__A1 (.I(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__B (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__I (.I(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05783__I (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__A1 (.I(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__I (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__I (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__I (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__A1 (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__A1 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__A1 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__A2 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__A1 (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A1 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A2 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__A1 (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__B (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__B1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05808__I (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__A2 (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__A1 (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__A1 (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__B1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__C1 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__A1 (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__A3 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A1 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__B1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__A3 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__A1 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__B1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__A2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__B1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__C1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05827__B (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__A2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__B1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A2 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__A1 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__A2 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05836__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05836__A2 (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__A1 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__A2 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__B (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__I (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__I (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__A2 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__A2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__I (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05853__A2 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A2 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__A2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__B2 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__A1 (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__A2 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__I (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__I (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A3 (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__I (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__A1 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__A2 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__A1 (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__A3 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__A2 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__I (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__I (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__A2 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A1 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A2 (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A2 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A3 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__A2 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__A1 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__A2 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__I (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A3 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__A1 (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__B1 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__I (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__A1 (.I(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__A3 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__A1 (.I(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__I (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__A1 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__A2 (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__B2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__B3 (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__I (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__I (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__I (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__I (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__I (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__I (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__I (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A1 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A2 (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A3 (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__A1 (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__A2 (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A1 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A2 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__I (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__I (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__I (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__I (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A1 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A2 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__A2 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__A3 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__A3 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__I (.I(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A1 (.I(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A2 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A3 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A1 (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A2 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__I (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__I (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__A1 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__B (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__A2 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A1 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A2 (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A2 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__A2 (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__B (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__C (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__A1 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A1 (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A2 (.I(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__I (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__I (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__I (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__I (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A2 (.I(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__I (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__I (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__I (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__A2 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__I (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__A1 (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A2 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__I (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__I (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__A1 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A2 (.I(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__I (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__I (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__I (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__I (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__A1 (.I(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__A2 (.I(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__I (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__I (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__A1 (.I(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__I (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__I (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__I (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__A1 (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A1 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__I (.I(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__I (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__I (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__I (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__A1 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A2 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__A1 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__B (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A2 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__A1 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__A2 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__C (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__A1 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__A2 (.I(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__B (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__A4 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__I (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__I (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A1 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A3 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__I (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A2 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__I (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__I (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__I (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A1 (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A1 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A2 (.I(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__B (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A3 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__I (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__B (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__I (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__A2 (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__I (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__B (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__I (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__I (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A2 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__B1 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A2 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__I (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A2 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__B1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__A2 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__I0 (.I(\as2650.regs[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__I1 (.I(\as2650.regs[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__S (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__I (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__I0 (.I(\as2650.regs[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__I1 (.I(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__I (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__I (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__I0 (.I(\as2650.regs[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__I1 (.I(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__I0 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__I1 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__I0 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__I1 (.I(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__I0 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__I1 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__S (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__I (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__I (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__I0 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__I1 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__S (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I0 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I1 (.I(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__S (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__I (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__I (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__I (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__I (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__S (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I0 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I1 (.I(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__S (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__S (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__I (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I0 (.I(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I1 (.I(\as2650.regs[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__I0 (.I(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__I1 (.I(\as2650.regs[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__I0 (.I(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__I1 (.I(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__S (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__I (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__A1 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__I (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__A2 (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__A1 (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__A2 (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__A3 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__A4 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__I (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__A1 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A2 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__B (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A1 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A1 (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A2 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__A1 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__I (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A1 (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__I (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__I (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__A1 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__A2 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A1 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__I (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__I (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A1 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A2 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__I (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A3 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__B (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A1 (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__I (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A1 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__A2 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__I (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__A2 (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__I (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A2 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__A1 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A1 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__I (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__A2 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A2 (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A2 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A1 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A3 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__I (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__A2 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__B (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A2 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A2 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__B (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A1 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A1 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__I (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A1 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A2 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__I (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A2 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__B (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A1 (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__C (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A2 (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A2 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A1 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__B (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A2 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A2 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A1 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__I (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A1 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A2 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__A2 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A2 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A2 (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__A1 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A2 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__I (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A1 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A2 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__A1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A1 (.I(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__A1 (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__A2 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__I (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__B1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__B2 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A1 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__I (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__I (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__I (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__I (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__B2 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__I (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__I (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__I (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__I (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__I (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__B1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__B1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__I (.I(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__B1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__I (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__B2 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__I (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__A2 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__I (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__I (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__I (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__B2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A2 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__B2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A2 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__B2 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A2 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__I (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__B1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__C (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__I (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__I (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__I (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__I (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__B1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__C (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__I (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__B1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__C (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__B1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__C (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__I (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__B1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__I (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__I (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__I (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__B1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__B1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__I (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__B1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__I (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__I (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__I (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__I (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__I (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__I (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__I (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__I (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__I (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__I (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__I (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__I (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__I (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A3 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A3 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A3 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__I (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__I (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__I (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__I (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A2 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__C (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A2 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__I (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__I (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A2 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__I (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__I (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__A3 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__A1 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A4 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A1 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A2 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__A1 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__I (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A2 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__I (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__I (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__I (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__I (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__I (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__I (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__I (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__I (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__I (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__I (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__I (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A1 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__A1 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A1 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__A1 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__I (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__I (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__I (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__I (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A2 (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__B (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A2 (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__B (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__A2 (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__B (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__I (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__I (.I(\as2650.PC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A2 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A1 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A1 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A2 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A1 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__I (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__I (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__I (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__I (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A1 (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A2 (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A2 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A2 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__I (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A1 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__I (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__I (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__I (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__A1 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__A2 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__I (.I(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__I (.I(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A2 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A2 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__I (.I(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__I (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A2 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A1 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A2 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__I (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A2 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__I (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__I (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A2 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A1 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A2 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A1 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A2 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__A2 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__I (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A2 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__I (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(\as2650.PC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A2 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A3 (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A1 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__I (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A1 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A2 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__A2 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__I (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__I (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__I (.I(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A1 (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A2 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A2 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__I (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A1 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A2 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__I (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A1 (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A2 (.I(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A2 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A2 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__I (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__I (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A1 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A2 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__A2 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__I (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A1 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A2 (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__I (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__I (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A2 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__A2 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A2 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__I (.I(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A1 (.I(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A2 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__I (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A2 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__I (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__I (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A1 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__I (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__I0 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__I1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A1 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A2 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__I (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A1 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__I0 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__A1 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__I (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__A1 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__I (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A2 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A2 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A2 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__I (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__A1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A1 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__A2 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__I (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__A2 (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__I0 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A1 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A1 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A2 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A2 (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A1 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__I (.I(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A1 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__B (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__I (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__I (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A1 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A1 (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__B (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__I (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A1 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__A1 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__B (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__I (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A2 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__I (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A1 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A1 (.I(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__I (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__I (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A3 (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__I (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A2 (.I(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A2 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A1 (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A1 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A2 (.I(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__B (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A2 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__S (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A2 (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A2 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A2 (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A3 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__I (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__I (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A2 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__I (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__I (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A1 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__I (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__A2 (.I(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A2 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A1 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__I (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A1 (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__I0 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A1 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__B2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__B (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__C (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A1 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A2 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A1 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A1 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__I (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A2 (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A2 (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__I (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__I (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__I (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07056__I (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__A1 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A3 (.I(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__A3 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__I (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A1 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A3 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A3 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__B (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A1 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A3 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A1 (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__I (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A2 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A3 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07077__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__A1 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A2 (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A3 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__A1 (.I(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__A2 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A2 (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__I (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__I (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__I (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__A2 (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A1 (.I(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A2 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A2 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A3 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A1 (.I(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A2 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__I (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A2 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__B (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A1 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A1 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__I (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__I (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A1 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A2 (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A2 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__A2 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__B (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__A1 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__C (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__I (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A1 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__A1 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__I (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__I (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__I (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A1 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__I (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__I (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__A2 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__B1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__B2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__A2 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__I (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__I (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__A1 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A1 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A2 (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A1 (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A2 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__B (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__C (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A2 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A1 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A2 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__I (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A2 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__B1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__B2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A2 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__I (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A2 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__I0 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__I1 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A2 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__I0 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__I1 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__S (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__C (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A1 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A1 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__C (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__I (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A2 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__B (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A1 (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__A1 (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A1 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__A2 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A1 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__I (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__I (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A2 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__B1 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__B2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__I (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A2 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__C (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A1 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__I (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__I0 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__I1 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__B2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A1 (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A2 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A2 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A3 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__A1 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A1 (.I(\as2650.regs[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A2 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__B1 (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__B2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__A2 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__I (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__I (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A2 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I0 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__S (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__I0 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__I1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__S (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A1 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A1 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__A1 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__I (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__A1 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__B2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__A1 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__A2 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A1 (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__I (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A1 (.I(\as2650.regs[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__B1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A2 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__A1 (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__A2 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__I0 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__I1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__S (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__I0 (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__I1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__S (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A1 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__A1 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__C (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A1 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A1 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A1 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A1 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__A2 (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__A1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__A2 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__I (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__A1 (.I(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__A2 (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__I (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__I (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A2 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A1 (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A2 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__A2 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A1 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__C (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A1 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__A1 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A1 (.I(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A2 (.I(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__B (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A2 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__B (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A1 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__C (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A1 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A2 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__I0 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__S (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__A1 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__A2 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__I (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__I (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__B1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A2 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__I (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__I (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__I (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A2 (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__A2 (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A2 (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A2 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__I (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A2 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A2 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A2 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A2 (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__A2 (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A2 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A2 (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A2 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A1 (.I(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A2 (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A2 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A2 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A2 (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A1 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__I (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__I (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__I (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A2 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A2 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A2 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__A1 (.I(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A2 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A1 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A1 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__I (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__A3 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__I (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__I (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__I (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__A2 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__A2 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A2 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__I (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A2 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A2 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A2 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A1 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A1 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__I (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__I (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__I (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__I (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__I (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A2 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A2 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__I (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A2 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__I (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A2 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__I (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A2 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__I (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A2 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__I (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A2 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__I (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__I (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__I (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__I (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__I (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A1 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A2 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__I (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__A1 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A1 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A2 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__I (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__I (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__I (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A3 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__I (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__I (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__I (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A2 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A2 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A2 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A2 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__I (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A2 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A2 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A2 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A2 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__A1 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A2 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A1 (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__B (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A1 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__B (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A1 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__B (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__I (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A1 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A1 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__A2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A2 (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A1 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A2 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__B (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A1 (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__I (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A1 (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A2 (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A1 (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A3 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A4 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__B1 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A1 (.I(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A2 (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__B (.I(\as2650.instruction_args_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A2 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__I (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A1 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A3 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__I (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__I (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__I (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__B (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__I (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__B1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A2 (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__B (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A3 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__I0 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__I1 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A2 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A3 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A1 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A2 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__I (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__I0 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__I1 (.I(\as2650.instruction_args_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A1 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__B (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A1 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A2 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__B1 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__I0 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__I1 (.I(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__S (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__I0 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__I1 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__B2 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__I (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A1 (.I(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__B1 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__C (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A1 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__I0 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__I1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A2 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__A2 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__I (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A1 (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A2 (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A3 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__A2 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A1 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A2 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A2 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__I (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__B1 (.I(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A1 (.I(\as2650.instruction_args_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__B1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__I0 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__I1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__I (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A1 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A2 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A2 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A1 (.I(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A1 (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__B1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__B2 (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__I (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__C (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__I (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A2 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__I (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__I (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__I0 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__I1 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__I (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A2 (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__B (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A1 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__B1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__B2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A2 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__I (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__I (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A2 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__B1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__B (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__A2 (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A2 (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__B (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A1 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__B1 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__I (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A2 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A1 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__B2 (.I(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A2 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__B1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__B2 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A1 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__I (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__I (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__I (.I(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A1 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__I (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__B1 (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__B1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__B2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A1 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__I (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__B1 (.I(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__B1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__B2 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A1 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__I (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__B (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A2 (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__B1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__B2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A1 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__I0 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__I1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__S (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__B2 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A1 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A1 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__A1 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__I (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__B2 (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A1 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A1 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__B (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A2 (.I(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A1 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__B (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__I (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__B (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__B2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A1 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__B2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__A1 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A2 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A1 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A1 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__I (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A1 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__C (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__B (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__I (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__I (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__I (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__B2 (.I(\as2650.instruction_args_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__I (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__B2 (.I(\as2650.instruction_args_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__I (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__I (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__B2 (.I(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__I (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__B2 (.I(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__I (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__B2 (.I(\as2650.instruction_args_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__B2 (.I(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__I (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__I (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__I (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__B1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A1 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__I (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__I (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__B1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__B2 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__B1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A1 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A1 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__B1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__B2 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A1 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A1 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A1 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__I (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A1 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A2 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A2 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A2 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A2 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A2 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A2 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A2 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A2 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A3 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A2 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__B (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A1 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__A2 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A2 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A3 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A4 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A2 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__I (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__I (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__I (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__I (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__I (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__I (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__I (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A2 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__B1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A2 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__I (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__I (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__I (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__I (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A2 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__B1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A1 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A1 (.I(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A2 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__B1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__B2 (.I(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__C (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__I (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__I (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A2 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__I0 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__I1 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A2 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__I (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__C (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A1 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A2 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A3 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A1 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__I (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A3 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__I (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A1 (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A3 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__I (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A1 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__B1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__B1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__C (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__B2 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__C (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A1 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A1 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A1 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__I (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__I (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__I (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__I (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__I (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__I (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__I (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__B1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__I (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__I (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__B1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A2 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__B1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A1 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A3 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A2 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__B1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__I (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__I (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__I (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__B1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__C (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A2 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__B1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__I (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__I (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__I (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__B1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__C (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__B1 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A2 (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__I0 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__I1 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__C (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__I (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__I (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__I (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__I (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__I (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__I (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A1 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__I (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__I (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__I (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__I (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__I (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__I (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A2 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A2 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__B (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A2 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A1 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__B (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A2 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A2 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A1 (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A2 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__B (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__I (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__I (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__I (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__I (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__I (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__I (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A2 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__I (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A2 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__B1 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__B1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A1 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__I (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__B1 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__B1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A1 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__I (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__I (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__I (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__I (.I(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A2 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__B1 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__C (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A2 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__B1 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__C (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__B1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A2 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A2 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__C (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A1 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__I (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A1 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__I (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__I (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__B (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__B2 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__I (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A1 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A3 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A2 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A3 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__B (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A1 (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__B2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__C (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__I (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__I (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A2 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A1 (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A3 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__B (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__I (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A2 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__B (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__I (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A2 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__B1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__I (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__I (.I(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A2 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__B1 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__B1 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A2 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__B1 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A1 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__B1 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__B1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__C (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__B1 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__B1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__C (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A2 (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__B (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A2 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A1 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__B (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__C (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A1 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__I (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__B1 (.I(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__B (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A1 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A2 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__I (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A1 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A2 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__I (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__I (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__I (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__B1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A2 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__B1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__I (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__I (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__B1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A2 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__B1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A2 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__B1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__I (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__B1 (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__C (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__A2 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__B1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__B2 (.I(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__C (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__B1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A2 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A2 (.I(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A2 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A1 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A2 (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__B2 (.I(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A2 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__B2 (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__B (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A2 (.I(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__I (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__I (.I(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__I (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__I (.I(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A2 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__B1 (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__C (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A2 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__B1 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__C (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__B1 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A2 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A2 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__I (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A1 (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A3 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A2 (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A1 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A1 (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__C (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A3 (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A1 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__B (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A2 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A2 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A2 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__B1 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__B1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A1 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__B1 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__B1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A1 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__B2 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__B1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__C (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A2 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__B1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__C (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__B1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A2 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A2 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A2 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A1 (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__A1 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__A2 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A2 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A1 (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__A1 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__B2 (.I(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__B2 (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__I (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__B (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__I (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__B1 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A2 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__B1 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__B1 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__B1 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__I (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__I (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__I (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__C (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A2 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__B1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__C (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A1 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__B1 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__A2 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__A2 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__I (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__I (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__A2 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A1 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__B (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A1 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A2 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__A1 (.I(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A2 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A2 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__I (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__A2 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A1 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A1 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__B (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A1 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__B (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A1 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__B2 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__B1 (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A1 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__A2 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__B2 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__B1 (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__B2 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__A1 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A1 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__B1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__B2 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__I (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__B1 (.I(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__C (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__B1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__B1 (.I(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__B2 (.I(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__C (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A1 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__C (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A2 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A1 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A2 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A3 (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__B (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A1 (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A2 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A2 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__C (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A1 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__B1 (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__B (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A1 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A2 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__B1 (.I(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A2 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__B1 (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A2 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__B1 (.I(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A2 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__B1 (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__A2 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__B1 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__C (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__B1 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__C (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A2 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__B (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A2 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__C (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__B1 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__B (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__B1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__A2 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__B1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A1 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__B1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__B1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__B1 (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A1 (.I(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A2 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__B1 (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__C (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__B1 (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__A2 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__B1 (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__C (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__I (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A1 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A2 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A2 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A1 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A2 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A2 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__B (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__B2 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A2 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__B2 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__C (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__I (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__B (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A2 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A1 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__I (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__I (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__I (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__B1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__B1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__B1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__I (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__B1 (.I(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A1 (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__B1 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__I (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__C (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__B1 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__C (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A2 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A2 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__B (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A1 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A2 (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__B2 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__I0 (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__S (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A1 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__B2 (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__C (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A1 (.I(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__B1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__B2 (.I(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__B1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__B1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__B1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A1 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__B1 (.I(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__B1 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__C (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__B1 (.I(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A2 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__B1 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__C (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__I0 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__I1 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A2 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A2 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A1 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A2 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A2 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A2 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__C (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A3 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__B2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__B (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A1 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__I (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__B1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__B1 (.I(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A2 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__B1 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A2 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__B1 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A1 (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__B1 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__C (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__C (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__B1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A2 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__B2 (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__C (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__B2 (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__B (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A2 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__B1 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A2 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__B1 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A2 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__B1 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A2 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__B1 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__C (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__C (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__B1 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A2 (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__C (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A1 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__B (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__B2 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__B (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A1 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__B1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__I (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A1 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__I (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A2 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A3 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A2 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__A2 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A2 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A1 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A4 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A2 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A3 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A4 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__C (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__I (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__I (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__I (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A2 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A3 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A2 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A1 (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A2 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__B (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A2 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A1 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A2 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A4 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A2 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A3 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A2 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__I (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A1 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A2 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__B (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__B (.I(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__C (.I(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A1 (.I(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A2 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__C (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A1 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A3 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__I (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A2 (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__B (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__I (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__B2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__I (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__I (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A2 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A2 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__I (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__I (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A2 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A2 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A1 (.I(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A2 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__C (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__B2 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A1 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A1 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__B (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__B2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__B2 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A1 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__B (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__B2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A1 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A1 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A2 (.I(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A2 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A1 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A2 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A1 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A1 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A1 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A2 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__I1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__B2 (.I(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__C (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A2 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A3 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A1 (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A2 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A2 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A2 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__B1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A2 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__B1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__B2 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A1 (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A2 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__B1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A2 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__B1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A1 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A2 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A2 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A1 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A2 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A2 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__B1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__B2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A2 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A3 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A3 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__B2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A2 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A3 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A1 (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A4 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A1 (.I(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A2 (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A1 (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A1 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A3 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A4 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A2 (.I(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A2 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A1 (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A1 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A3 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A4 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__B (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A2 (.I(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A2 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__B1 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__B2 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A2 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A1 (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A2 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__B1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__B2 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A2 (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__B1 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__B2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__B1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__C1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__C2 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A2 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A3 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__B2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A1 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A3 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A2 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A2 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A3 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A1 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A1 (.I(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A1 (.I(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A1 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A3 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A4 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A1 (.I(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A2 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__B1 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__B2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A1 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A1 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A2 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A1 (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A2 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A2 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A2 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A3 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A4 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__I (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A2 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A2 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A1 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A2 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A1 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A4 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A1 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A2 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A1 (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A2 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A3 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A4 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A2 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__B2 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A1 (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A2 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A2 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__B1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A2 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A1 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__A1 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A2 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A2 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__I (.I(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__B1 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A1 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A2 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A1 (.I(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A1 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__B2 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A2 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A1 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A2 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A1 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A2 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__B2 (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__A3 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A3 (.I(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A3 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A1 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__B1 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__C2 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__B1 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__B2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A1 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__B1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__C (.I(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__I (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A1 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A2 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__A1 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A2 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A1 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A2 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A2 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__C (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__B (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A1 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__C (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__B (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A1 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A2 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A3 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A4 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A3 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__C (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A1 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A3 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A1 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__B1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A1 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__B (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A1 (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A2 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__I (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A2 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__B (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__B (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A1 (.I(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A2 (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__C (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A2 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__I (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A2 (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__I (.I(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A1 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__I (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__I (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A1 (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A2 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A3 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__B (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A1 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A2 (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__B (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__B1 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__B2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__C (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A2 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__I (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__I (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A1 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A3 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A1 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__B1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__B2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A2 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__C (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A2 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__A1 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A2 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__B2 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A1 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__C (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A2 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__B2 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A1 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__C (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__B (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__B2 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A1 (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A2 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__B2 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__B2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__B2 (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A2 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A1 (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A1 (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__A1 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__B2 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A2 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__C (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__A1 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__B2 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__B (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A2 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__B (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__C (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A2 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__I (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__I (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__I (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A2 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A2 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A1 (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A3 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__I (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A2 (.I(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A1 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A2 (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A2 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A2 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A3 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A1 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A2 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__B1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__B2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A1 (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A2 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A2 (.I(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A2 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A1 (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A1 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__C (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A2 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A1 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__B1 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__B2 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__I (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__I (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A1 (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A1 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A2 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A1 (.I(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__I (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__B1 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__B2 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A1 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__I (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__I (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A2 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A1 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A1 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__B1 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__B2 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__I (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__A1 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A2 (.I(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A1 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A1 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__B1 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__B2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__A1 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A2 (.I(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A1 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__B1 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__B2 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__I (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A1 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A1 (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A1 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__B1 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__B2 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A1 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A1 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A1 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A2 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A1 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A2 (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A1 (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A3 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__I (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A1 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A2 (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__I (.I(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__I (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A1 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A2 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__B (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__I (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A1 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__A1 (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A1 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A1 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__I (.I(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__I (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__I (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A1 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__A1 (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__I (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__A1 (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__B2 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A2 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A2 (.I(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__I (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__A2 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__B2 (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A1 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A2 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A1 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__B2 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A2 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__B1 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A1 (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__B2 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__A1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__B (.I(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A1 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__B1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__B2 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__B1 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__B2 (.I(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__A1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__B1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__B2 (.I(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__A1 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A2 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__B1 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A1 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__B2 (.I(\as2650.regs[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A1 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A2 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A1 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__B1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__B2 (.I(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A1 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A1 (.I(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A3 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__B2 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A1 (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__B2 (.I(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A1 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A2 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__A1 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__B2 (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__I (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A2 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A1 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__B2 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__B2 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A1 (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__B2 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__B2 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__B2 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A1 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__B2 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__A1 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__B2 (.I(\as2650.regs[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__B2 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__B2 (.I(\as2650.regs[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__B2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A1 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__B2 (.I(\as2650.regs[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__B2 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__B2 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__I (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A1 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A1 (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__I1 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A2 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A3 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A2 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__B (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A1 (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__I (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A1 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__B2 (.I(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A2 (.I(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__B2 (.I(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A1 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A2 (.I(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__B2 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A1 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A1 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A2 (.I(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__B2 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__A1 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A1 (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A2 (.I(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__B2 (.I(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A1 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A1 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__B2 (.I(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A1 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A1 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__A1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A2 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A1 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__I0 (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__I0 (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A2 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A3 (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__I (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A3 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A4 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__I (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A2 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__B (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__I (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A1 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__A1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__A1 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A1 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__I (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__I (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__I (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A1 (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__B2 (.I(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__B2 (.I(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__A1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__B2 (.I(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A1 (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A1 (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A2 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A2 (.I(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__A2 (.I(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__A1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A2 (.I(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__A2 (.I(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__A2 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__A2 (.I(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A2 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A2 (.I(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A2 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A2 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__A2 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__I (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A2 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__I (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__I (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__I (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__I (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A1 (.I(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__I (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A1 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__I (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__I (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__I (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A1 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A1 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__I (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A1 (.I(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__I (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A1 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__I (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__I (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__I (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A2 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A2 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__I (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A2 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A1 (.I(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A2 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__I (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A2 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A2 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__I (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A2 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A2 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__I (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__I (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__I (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__I (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__I (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A2 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__I (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A2 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A2 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A2 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A1 (.I(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A2 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__I (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A1 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A1 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A1 (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A1 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__I (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A2 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A2 (.I(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A2 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A1 (.I(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A2 (.I(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A2 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A2 (.I(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A2 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A2 (.I(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__I (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__I (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__I (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__I (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__I (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A1 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__A1 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A1 (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__A1 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__I (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__I (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A1 (.I(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__I (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__I (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__I (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A1 (.I(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A1 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__I (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A1 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__I (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A1 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A2 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__C (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__I (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A1 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A2 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__I (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A1 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A2 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__B (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__I (.I(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A1 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A1 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A1 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__I (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__I (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__I (.I(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A1 (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A1 (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__B2 (.I(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__I (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__I (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A1 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__I (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__I (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A1 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__A1 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A1 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A1 (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A1 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__I (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__I (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A1 (.I(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__I (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__I (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A1 (.I(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A1 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__I (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A3 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__I (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__I (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__I (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A2 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__I (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A2 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__I (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A2 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__I (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A2 (.I(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__I (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__I (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A2 (.I(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A1 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A2 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__A2 (.I(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A1 (.I(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A2 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__I (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A2 (.I(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A2 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__I (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A2 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__I (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A1 (.I(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__I (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__I (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__I (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A2 (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A1 (.I(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A2 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__I (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A1 (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__I (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A1 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A1 (.I(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__I (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__A1 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__I (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__A1 (.I(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A1 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A1 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__A1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A1 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__I (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A1 (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A1 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__I (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A1 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A1 (.I(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__A1 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__A1 (.I(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__A2 (.I(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A2 (.I(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A2 (.I(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A2 (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A1 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A2 (.I(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__A2 (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A1 (.I(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A2 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__A2 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__I (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__I (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__A1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A1 (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__A1 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__I (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__I (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A1 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A1 (.I(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__I (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__I (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A1 (.I(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__A1 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__I (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__I (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__A1 (.I(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A1 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A1 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__D (.I(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__D (.I(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__CLK (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__D (.I(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__D (.I(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__D (.I(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__D (.I(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__D (.I(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__D (.I(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__D (.I(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__D (.I(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__CLK (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__CLK (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__CLK (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__CLK (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__CLK (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold102_I (.I(wbs_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold106_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold113_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold116_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold119_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold122_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold125_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold128_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold131_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold134_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold137_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold140_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold143_I (.I(wbs_adr_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold144_I (.I(wbs_adr_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold148_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold150_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold151_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold152_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold153_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold32_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold36_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold40_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold44_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold48_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold52_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold56_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold60_I (.I(wbs_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold64_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold68_I (.I(wbs_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold72_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold79_I (.I(wbs_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold83_I (.I(wbs_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold87_I (.I(wbs_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold91_I (.I(wbs_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold95_I (.I(wbs_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output74_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output84_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output89_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output90_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output91_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer17_I (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer21_I (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer25_I (.I(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer27_I (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer29_I (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer5_I (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer8_I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_510 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05231_ (.I(net11),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05232_ (.A1(_00502_),
    .A2(net1),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _05233_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(_00503_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05234_ (.I(_00504_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05235_ (.I(_00505_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05236_ (.I(_00506_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05237_ (.I(_00507_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05238_ (.I(_00508_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05239_ (.I(_00509_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05240_ (.I(\as2650.cycle[3] ),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05241_ (.I(_00511_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05242_ (.I(\as2650.cycle[0] ),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05243_ (.I(_00513_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05244_ (.I(_00514_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05245_ (.I(_00515_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05246_ (.I(_00516_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _05247_ (.I(net8),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05248_ (.A1(_00518_),
    .A2(_00516_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05249_ (.A1(\as2650.insin[2] ),
    .A2(_00517_),
    .B(_00519_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05250_ (.I(_00520_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05251_ (.I(\as2650.extend ),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05252_ (.I(_00522_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05253_ (.I(_00523_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05254_ (.I(\as2650.indirect_cyc ),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05255_ (.I(_00525_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05256_ (.A1(_00524_),
    .A2(_00526_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05257_ (.I(_00527_),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05258_ (.I(net4),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05259_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(_00503_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05260_ (.I(\as2650.cycle[5] ),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05261_ (.I(_00531_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05262_ (.I(_00532_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05263_ (.I(_00533_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05264_ (.I(_00534_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05265_ (.I(\as2650.instruction_args_latch[13] ),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05266_ (.A1(_00523_),
    .A2(_00526_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05267_ (.A1(_00536_),
    .A2(_00537_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05268_ (.A1(\as2650.page_reg[0] ),
    .A2(_00527_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05269_ (.A1(_00535_),
    .A2(_00538_),
    .A3(_00539_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05270_ (.I(\as2650.relative_cyc ),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05271_ (.A1(_00541_),
    .A2(_00525_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05272_ (.I(_00542_),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05273_ (.I(_00514_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05274_ (.A1(_00544_),
    .A2(\as2650.cycle[3] ),
    .A3(\as2650.cycle[2] ),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05275_ (.I(_00545_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05276_ (.A1(\as2650.relative_cyc ),
    .A2(\as2650.indirect_cyc ),
    .A3(\as2650.cycle[5] ),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05277_ (.I(_00547_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05278_ (.A1(_00546_),
    .A2(_00548_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05279_ (.I(_00549_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05280_ (.A1(\as2650.indirect_target[7] ),
    .A2(_00543_),
    .B1(_00550_),
    .B2(\as2650.PC[7] ),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05281_ (.I(\as2650.indirect_target[6] ),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05282_ (.A1(\as2650.relative_cyc ),
    .A2(\as2650.indirect_cyc ),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05283_ (.I(_00553_),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05284_ (.A1(_00545_),
    .A2(_00547_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05285_ (.I(_00555_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _05286_ (.I(\as2650.PC[6] ),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _05287_ (.A1(_00552_),
    .A2(_00554_),
    .B1(_00556_),
    .B2(_00557_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05288_ (.I(\as2650.indirect_target[5] ),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _05289_ (.I(\as2650.PC[5] ),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _05290_ (.A1(_00559_),
    .A2(_00554_),
    .B1(_00556_),
    .B2(_00560_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05291_ (.I(\as2650.PC[3] ),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05292_ (.I(\as2650.indirect_target[3] ),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _05293_ (.A1(_00562_),
    .A2(_00545_),
    .A3(_00548_),
    .B1(_00553_),
    .B2(_00563_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05294_ (.I(\as2650.cycle[2] ),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _05295_ (.I(_00565_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05296_ (.A1(\as2650.relative_cyc ),
    .A2(\as2650.indirect_cyc ),
    .A3(_00531_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05297_ (.A1(_00541_),
    .A2(_00525_),
    .B(\as2650.indirect_target[1] ),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05298_ (.A1(_00541_),
    .A2(_00525_),
    .B(\as2650.indirect_target[0] ),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05299_ (.A1(_00566_),
    .A2(_00567_),
    .A3(_00568_),
    .A4(_00569_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _05300_ (.I(\as2650.PC[2] ),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05301_ (.I(\as2650.indirect_target[2] ),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _05302_ (.A1(_00571_),
    .A2(_00546_),
    .A3(_00548_),
    .B1(_00554_),
    .B2(_00572_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05303_ (.A1(_00564_),
    .A2(_00570_),
    .A3(_00573_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05304_ (.I(\as2650.PC[4] ),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05305_ (.A1(\as2650.indirect_target[4] ),
    .A2(_00542_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05306_ (.A1(_00575_),
    .A2(_00555_),
    .B(_00576_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05307_ (.A1(_00574_),
    .A2(_00577_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _05308_ (.A1(_00558_),
    .A2(_00561_),
    .A3(_00578_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05309_ (.A1(\as2650.indirect_target[8] ),
    .A2(_00543_),
    .B1(_00550_),
    .B2(\as2650.PC[8] ),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05310_ (.A1(_00551_),
    .A2(_00579_),
    .A3(_00580_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05311_ (.I(_00543_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05312_ (.A1(\as2650.indirect_target[9] ),
    .A2(_00582_),
    .B1(_00550_),
    .B2(\as2650.PC[9] ),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05313_ (.I(_00583_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05314_ (.A1(_00581_),
    .A2(_00584_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05315_ (.I(_00550_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05316_ (.A1(\as2650.indirect_target[10] ),
    .A2(_00582_),
    .B1(_00586_),
    .B2(\as2650.PC[10] ),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05317_ (.A1(\as2650.indirect_target[11] ),
    .A2(_00582_),
    .B1(_00586_),
    .B2(\as2650.PC[11] ),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05318_ (.A1(_00585_),
    .A2(_00587_),
    .A3(_00588_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05319_ (.I(_00582_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05320_ (.A1(\as2650.indirect_target[12] ),
    .A2(_00590_),
    .B1(_00586_),
    .B2(\as2650.PC[12] ),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05321_ (.I(_00591_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05322_ (.A1(_00589_),
    .A2(_00592_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05323_ (.I(_00586_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05324_ (.A1(\as2650.indirect_target[13] ),
    .A2(_00590_),
    .B1(_00594_),
    .B2(\as2650.page_reg[0] ),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05325_ (.A1(_00593_),
    .A2(_00595_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05326_ (.A1(_00593_),
    .A2(_00595_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05327_ (.I(_00531_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05328_ (.I(_00598_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05329_ (.A1(_00596_),
    .A2(_00597_),
    .B(_00599_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05330_ (.A1(_00540_),
    .A2(_00600_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05331_ (.I0(\as2650.insin[3] ),
    .I1(net9),
    .S(_00515_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05332_ (.I0(\as2650.insin[2] ),
    .I1(net8),
    .S(_00515_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05333_ (.A1(_00602_),
    .A2(_00603_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05334_ (.A1(_00526_),
    .A2(_00604_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _05335_ (.I(\as2650.extend ),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05336_ (.I0(\as2650.insin[4] ),
    .I1(net10),
    .S(_00544_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05337_ (.I0(\as2650.insin[5] ),
    .I1(net2),
    .S(_00515_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _05338_ (.A1(_00607_),
    .A2(_00608_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05339_ (.I0(\as2650.insin[7] ),
    .I1(net4),
    .S(_00544_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05340_ (.I0(\as2650.insin[6] ),
    .I1(net3),
    .S(_00544_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05341_ (.A1(_00610_),
    .A2(_00611_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05342_ (.I(_00607_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _05343_ (.A1(_00613_),
    .A2(_00602_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05344_ (.A1(\as2650.instruction_args_latch[13] ),
    .A2(\as2650.instruction_args_latch[14] ),
    .B(_00606_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _05345_ (.A1(_00606_),
    .A2(_00609_),
    .A3(_00612_),
    .B1(_00614_),
    .B2(_00615_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05346_ (.I(\as2650.indexed_cyc[1] ),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05347_ (.I(\as2650.indexed_cyc[0] ),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05348_ (.A1(_00605_),
    .A2(_00616_),
    .B(_00617_),
    .C(_00618_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05349_ (.A1(_00598_),
    .A2(_00619_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05350_ (.I(_00620_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05351_ (.I(_00541_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05352_ (.A1(_00622_),
    .A2(_00605_),
    .A3(_00616_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05353_ (.A1(_00621_),
    .A2(_00623_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05354_ (.I(_00624_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05355_ (.I(\as2650.indexed_cyc[1] ),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05356_ (.A1(_00626_),
    .A2(_00536_),
    .B(_00618_),
    .C(_00522_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05357_ (.I(\as2650.indexed_cyc[0] ),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05358_ (.I(\as2650.instruction_args_latch[14] ),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05359_ (.A1(_00628_),
    .A2(_00629_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05360_ (.A1(_00523_),
    .A2(_00617_),
    .A3(_00627_),
    .A4(_00630_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05361_ (.I(_00631_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05362_ (.A1(_00626_),
    .A2(\as2650.instruction_args_latch[13] ),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05363_ (.A1(_00628_),
    .A2(\as2650.instruction_args_latch[14] ),
    .B(\as2650.extend ),
    .C(_00617_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05364_ (.A1(_00522_),
    .A2(_00618_),
    .A3(_00633_),
    .A4(_00634_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05365_ (.I(_00635_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05366_ (.I(_00636_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05367_ (.I0(\as2650.insin[1] ),
    .I1(net7),
    .S(_00513_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _05368_ (.I(net242),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05369_ (.I0(\as2650.insin[0] ),
    .I1(net6),
    .S(\as2650.cycle[0] ),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05370_ (.I(_00640_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05371_ (.A1(_00641_),
    .A2(_00639_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05372_ (.I(_00642_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05373_ (.I(_00643_),
    .Z(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05374_ (.I(_00644_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05375_ (.I(\as2650.debug_psl[4] ),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05376_ (.I(_00646_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05377_ (.I(_00647_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05378_ (.I(_00648_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05379_ (.I(_00649_),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05380_ (.A1(\as2650.regs[3][7] ),
    .A2(_00645_),
    .B(_00650_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _05381_ (.A1(net239),
    .A2(_00641_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _05382_ (.I(_00652_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05383_ (.I(_00653_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05384_ (.I(\as2650.insin[0] ),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05385_ (.A1(net6),
    .A2(_00513_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _05386_ (.A1(_00655_),
    .A2(_00514_),
    .B(net240),
    .C(_00656_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05387_ (.I(_00657_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05388_ (.I(_00658_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05389_ (.I(_00659_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05390_ (.I(\as2650.insin[1] ),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05391_ (.A1(net7),
    .A2(_00513_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _05392_ (.A1(_00661_),
    .A2(_00514_),
    .B(_00662_),
    .C(_00640_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05393_ (.I(_00663_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05394_ (.I(_00664_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05395_ (.I(_00665_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _05396_ (.A1(\as2650.regs[0][7] ),
    .A2(_00654_),
    .B1(_00660_),
    .B2(\as2650.regs[2][7] ),
    .C1(_00666_),
    .C2(\as2650.regs[1][7] ),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05397_ (.A1(_00651_),
    .A2(_00667_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05398_ (.I(\as2650.regs[4][7] ),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05399_ (.A1(_00639_),
    .A2(_00641_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05400_ (.I(_00646_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05401_ (.I(_00671_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05402_ (.A1(\as2650.regs[7][7] ),
    .A2(_00644_),
    .B(_00672_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05403_ (.A1(\as2650.regs[6][7] ),
    .A2(_00660_),
    .B1(_00666_),
    .B2(\as2650.regs[5][7] ),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05404_ (.A1(_00669_),
    .A2(_00670_),
    .B(_00673_),
    .C(_00674_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05405_ (.A1(_00668_),
    .A2(_00675_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05406_ (.I(_00646_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05407_ (.A1(\as2650.regs[1][1] ),
    .A2(_00665_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05408_ (.I(_00657_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05409_ (.A1(\as2650.regs[2][1] ),
    .A2(_00679_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _05410_ (.I(_00642_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _05411_ (.I(_00652_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _05412_ (.A1(\as2650.regs[3][1] ),
    .A2(_00681_),
    .B1(_00682_),
    .B2(\as2650.regs[0][1] ),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05413_ (.A1(_00677_),
    .A2(_00678_),
    .A3(_00680_),
    .A4(_00683_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05414_ (.I(\as2650.debug_psl[4] ),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05415_ (.A1(\as2650.regs[7][1] ),
    .A2(_00681_),
    .B(_00685_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05416_ (.I(_00663_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05417_ (.A1(\as2650.regs[5][1] ),
    .A2(_00687_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05418_ (.A1(\as2650.regs[6][1] ),
    .A2(_00679_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05419_ (.A1(\as2650.regs[4][1] ),
    .A2(_00682_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05420_ (.A1(_00686_),
    .A2(_00688_),
    .A3(_00689_),
    .A4(_00690_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05421_ (.A1(_00684_),
    .A2(_00691_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05422_ (.A1(\as2650.regs[1][0] ),
    .A2(_00664_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05423_ (.A1(\as2650.regs[2][0] ),
    .A2(_00658_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _05424_ (.A1(\as2650.regs[3][0] ),
    .A2(_00642_),
    .B1(_00652_),
    .B2(\as2650.regs[0][0] ),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05425_ (.A1(_00677_),
    .A2(_00693_),
    .A3(_00694_),
    .A4(_00695_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05426_ (.A1(\as2650.regs[7][0] ),
    .A2(_00681_),
    .B(_00685_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05427_ (.A1(\as2650.regs[5][0] ),
    .A2(_00664_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05428_ (.A1(net385),
    .A2(\as2650.regs[6][0] ),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05429_ (.A1(_00682_),
    .A2(\as2650.regs[4][0] ),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05430_ (.A1(_00697_),
    .A2(_00698_),
    .A3(_00699_),
    .A4(_00700_),
    .Z(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05431_ (.A1(_00696_),
    .A2(net245),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05432_ (.A1(\as2650.regs[3][2] ),
    .A2(_00681_),
    .B(_00648_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _05433_ (.A1(\as2650.regs[0][2] ),
    .A2(_00682_),
    .B1(_00679_),
    .B2(\as2650.regs[2][2] ),
    .C1(_00687_),
    .C2(\as2650.regs[1][2] ),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05434_ (.A1(_00703_),
    .A2(_00704_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05435_ (.A1(\as2650.regs[7][2] ),
    .A2(_00643_),
    .B(_00685_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _05436_ (.A1(\as2650.regs[4][2] ),
    .A2(_00653_),
    .B1(_00679_),
    .B2(\as2650.regs[6][2] ),
    .C1(_00687_),
    .C2(\as2650.regs[5][2] ),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05437_ (.A1(_00706_),
    .A2(_00707_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05438_ (.A1(_00705_),
    .A2(net248),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05439_ (.I(_00647_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05440_ (.A1(\as2650.regs[3][3] ),
    .A2(_00643_),
    .B(_00710_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _05441_ (.A1(\as2650.regs[0][3] ),
    .A2(_00653_),
    .B1(_00659_),
    .B2(\as2650.regs[2][3] ),
    .C1(_00687_),
    .C2(\as2650.regs[1][3] ),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05442_ (.A1(_00712_),
    .A2(_00711_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05443_ (.A1(\as2650.regs[7][3] ),
    .A2(_00643_),
    .B(_00677_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _05444_ (.A1(\as2650.regs[4][3] ),
    .A2(_00653_),
    .B1(_00659_),
    .B2(\as2650.regs[6][3] ),
    .C1(_00665_),
    .C2(\as2650.regs[5][3] ),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05445_ (.A1(_00714_),
    .A2(_00715_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _05446_ (.A1(_00713_),
    .A2(_00716_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05447_ (.I(_00717_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05448_ (.A1(_00692_),
    .A2(_00702_),
    .A3(_00709_),
    .A4(_00718_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05449_ (.I(_00664_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05450_ (.A1(\as2650.regs[1][5] ),
    .A2(_00720_),
    .B(_00710_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05451_ (.I(_00652_),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05452_ (.I(_00658_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05453_ (.I(_00642_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _05454_ (.A1(\as2650.regs[0][5] ),
    .A2(_00722_),
    .B1(_00723_),
    .B2(\as2650.regs[2][5] ),
    .C1(\as2650.regs[3][5] ),
    .C2(_00724_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05455_ (.A1(_00721_),
    .A2(_00725_),
    .Z(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05456_ (.I(_00646_),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05457_ (.A1(\as2650.regs[5][5] ),
    .A2(_00720_),
    .B(_00727_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _05458_ (.A1(\as2650.regs[4][5] ),
    .A2(_00722_),
    .B1(_00723_),
    .B2(\as2650.regs[6][5] ),
    .C1(\as2650.regs[7][5] ),
    .C2(_00724_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05459_ (.A1(_00728_),
    .A2(_00729_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05460_ (.A1(_00726_),
    .A2(_00730_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05461_ (.I(_00731_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05462_ (.A1(\as2650.regs[1][4] ),
    .A2(_00665_),
    .B(_00710_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _05463_ (.A1(\as2650.regs[0][4] ),
    .A2(_00722_),
    .B1(_00659_),
    .B2(\as2650.regs[2][4] ),
    .C1(\as2650.regs[3][4] ),
    .C2(_00724_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05464_ (.A1(_00733_),
    .A2(_00734_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05465_ (.I(_00685_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05466_ (.A1(\as2650.regs[5][4] ),
    .A2(_00720_),
    .B(_00736_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _05467_ (.A1(\as2650.regs[4][4] ),
    .A2(_00722_),
    .B1(_00723_),
    .B2(\as2650.regs[6][4] ),
    .C1(\as2650.regs[7][4] ),
    .C2(_00724_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05468_ (.A1(_00737_),
    .A2(_00738_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05469_ (.A1(_00735_),
    .A2(_00739_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05470_ (.I(_00740_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05471_ (.A1(_00732_),
    .A2(_00741_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05472_ (.A1(\as2650.regs[1][6] ),
    .A2(_00720_),
    .B(_00649_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _05473_ (.A1(\as2650.regs[0][6] ),
    .A2(_00654_),
    .B1(_00723_),
    .B2(\as2650.regs[2][6] ),
    .C1(\as2650.regs[3][6] ),
    .C2(_00644_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05474_ (.A1(_00743_),
    .A2(_00744_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05475_ (.I(_00736_),
    .Z(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05476_ (.A1(\as2650.regs[5][6] ),
    .A2(_00666_),
    .B(_00746_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _05477_ (.A1(\as2650.regs[4][6] ),
    .A2(_00654_),
    .B1(_00660_),
    .B2(\as2650.regs[6][6] ),
    .C1(\as2650.regs[7][6] ),
    .C2(_00644_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05478_ (.A1(_00747_),
    .A2(_00748_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05479_ (.A1(_00745_),
    .A2(_00749_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05480_ (.A1(_00676_),
    .A2(net234),
    .A3(_00742_),
    .A4(_00750_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05481_ (.A1(_00727_),
    .A2(_00678_),
    .A3(_00680_),
    .A4(_00683_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05482_ (.A1(_00686_),
    .A2(_00688_),
    .A3(_00689_),
    .A4(_00690_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05483_ (.A1(_00753_),
    .A2(_00752_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05484_ (.I(_00754_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05485_ (.A1(_00746_),
    .A2(_00693_),
    .A3(_00694_),
    .A4(_00695_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05486_ (.A1(_00697_),
    .A2(_00698_),
    .A3(_00699_),
    .A4(net259),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05487_ (.A1(_00757_),
    .A2(_00756_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05488_ (.A1(_00705_),
    .A2(_00708_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05489_ (.A1(_00713_),
    .A2(_00716_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05490_ (.A1(_00755_),
    .A2(_00758_),
    .A3(_00759_),
    .A4(_00760_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05491_ (.I(_00761_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05492_ (.A1(_00726_),
    .A2(_00730_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05493_ (.A1(_00735_),
    .A2(_00739_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05494_ (.A1(_00764_),
    .A2(_00763_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05495_ (.A1(_00745_),
    .A2(_00749_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05496_ (.A1(_00668_),
    .A2(_00675_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05497_ (.A1(_00762_),
    .A2(_00765_),
    .A3(_00766_),
    .B(_00767_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _05498_ (.A1(_00637_),
    .A2(_00751_),
    .A3(_00768_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05499_ (.I(_00767_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05500_ (.A1(_00637_),
    .A2(_00770_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05501_ (.I(_00631_),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05502_ (.I(_00750_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05503_ (.I(_00718_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05504_ (.A1(_00684_),
    .A2(_00691_),
    .B1(_00696_),
    .B2(_00701_),
    .C1(_00705_),
    .C2(_00708_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05505_ (.I(_00775_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05506_ (.A1(_00774_),
    .A2(_00732_),
    .A3(_00741_),
    .A4(_00776_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05507_ (.A1(_00773_),
    .A2(_00777_),
    .B(_00676_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05508_ (.I(_00766_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _05509_ (.A1(_00717_),
    .A2(_00731_),
    .A3(_00740_),
    .A4(_00775_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05510_ (.A1(_00770_),
    .A2(_00779_),
    .A3(_00780_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05511_ (.A1(_00772_),
    .A2(_00778_),
    .A3(_00781_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05512_ (.A1(_00632_),
    .A2(_00769_),
    .A3(_00771_),
    .B(_00782_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05513_ (.I(_00531_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05514_ (.I(_00784_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05515_ (.A1(_00785_),
    .A2(\as2650.instruction_args_latch[7] ),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05516_ (.I(_00784_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05517_ (.A1(_00551_),
    .A2(_00579_),
    .B(_00787_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05518_ (.A1(_00551_),
    .A2(_00579_),
    .B(_00788_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05519_ (.A1(_00786_),
    .A2(_00789_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05520_ (.A1(_00625_),
    .A2(_00783_),
    .A3(_00790_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05521_ (.I(_00791_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05522_ (.A1(_00620_),
    .A2(_00623_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05523_ (.I(_00793_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05524_ (.I(_00676_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05525_ (.A1(_00637_),
    .A2(_00795_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05526_ (.A1(_00523_),
    .A2(_00617_),
    .A3(_00630_),
    .B(_00627_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05527_ (.I(_00797_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05528_ (.A1(_00751_),
    .A2(_00768_),
    .B(_00798_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05529_ (.A1(_00676_),
    .A2(_00779_),
    .A3(_00780_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05530_ (.A1(_00773_),
    .A2(_00777_),
    .B(_00770_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05531_ (.A1(_00632_),
    .A2(_00800_),
    .A3(_00801_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05532_ (.A1(_00632_),
    .A2(_00796_),
    .A3(_00799_),
    .B(_00802_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05533_ (.A1(_00786_),
    .A2(_00789_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05534_ (.A1(_00794_),
    .A2(_00803_),
    .B(_00804_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05535_ (.I(_00805_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05536_ (.A1(_00719_),
    .A2(_00742_),
    .B(_00766_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05537_ (.A1(_00761_),
    .A2(_00765_),
    .A3(_00750_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05538_ (.A1(_00797_),
    .A2(_00766_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05539_ (.A1(_00798_),
    .A2(_00807_),
    .A3(_00808_),
    .B(_00809_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05540_ (.A1(_00780_),
    .A2(_00750_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05541_ (.A1(_00811_),
    .A2(_00631_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _05542_ (.A1(_00772_),
    .A2(_00810_),
    .B(_00812_),
    .C(_00793_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05543_ (.A1(_00561_),
    .A2(_00578_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05544_ (.A1(_00558_),
    .A2(_00814_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05545_ (.A1(_00784_),
    .A2(\as2650.instruction_args_latch[6] ),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05546_ (.A1(_00599_),
    .A2(_00815_),
    .B(_00816_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05547_ (.A1(_00813_),
    .A2(_00817_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05548_ (.I(_00818_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05549_ (.A1(_00792_),
    .A2(_00806_),
    .A3(_00819_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05550_ (.A1(_00631_),
    .A2(_00636_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05551_ (.I(_00821_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05552_ (.A1(_00696_),
    .A2(net247),
    .B(_00822_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05553_ (.A1(_00696_),
    .A2(net246),
    .A3(_00821_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05554_ (.A1(_00824_),
    .A2(_00823_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05555_ (.I(\as2650.indirect_target[0] ),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05556_ (.A1(_00826_),
    .A2(_00566_),
    .A3(_00554_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05557_ (.I(_00548_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05558_ (.A1(\as2650.indirect_target[0] ),
    .A2(_00542_),
    .B1(_00828_),
    .B2(_00565_),
    .C1(_00549_),
    .C2(\as2650.PC[0] ),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05559_ (.A1(\as2650.instruction_args_latch[0] ),
    .A2(_00784_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05560_ (.A1(_00532_),
    .A2(_00827_),
    .A3(_00829_),
    .B(_00830_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05561_ (.A1(_00793_),
    .A2(_00825_),
    .A3(_00831_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05562_ (.A1(_00522_),
    .A2(_00618_),
    .A3(_00633_),
    .B(_00634_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05563_ (.A1(_00635_),
    .A2(_00756_),
    .A3(_00757_),
    .B(_00833_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _05564_ (.A1(_00754_),
    .A2(_00702_),
    .A3(_00834_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _05565_ (.A1(\as2650.indirect_target[1] ),
    .A2(_00543_),
    .B1(_00549_),
    .B2(\as2650.PC[1] ),
    .C(_00827_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05566_ (.A1(_00532_),
    .A2(\as2650.instruction_args_latch[1] ),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05567_ (.A1(_00532_),
    .A2(_00570_),
    .A3(_00836_),
    .B(_00837_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05568_ (.A1(_00794_),
    .A2(_00835_),
    .B(_00838_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05569_ (.I(_00835_),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05570_ (.A1(_00794_),
    .A2(_00840_),
    .A3(_00838_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05571_ (.A1(_00832_),
    .A2(_00839_),
    .B(_00841_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05572_ (.I(_00624_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05573_ (.I(_00758_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05574_ (.A1(_00755_),
    .A2(_00844_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05575_ (.I(_00709_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05576_ (.I(_00702_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05577_ (.A1(_00692_),
    .A2(_00847_),
    .A3(_00709_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05578_ (.A1(_00845_),
    .A2(_00846_),
    .B(_00848_),
    .C(_00798_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05579_ (.A1(_00752_),
    .A2(_00753_),
    .B1(_00756_),
    .B2(net260),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05580_ (.A1(_00759_),
    .A2(_00850_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05581_ (.A1(_00759_),
    .A2(_00822_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05582_ (.A1(_00833_),
    .A2(_00851_),
    .B(_00852_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05583_ (.A1(_00570_),
    .A2(_00573_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05584_ (.A1(_00570_),
    .A2(_00573_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05585_ (.A1(_00787_),
    .A2(_00855_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05586_ (.A1(_00785_),
    .A2(\as2650.instruction_args_latch[2] ),
    .B1(_00854_),
    .B2(_00856_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05587_ (.A1(_00843_),
    .A2(_00849_),
    .A3(_00853_),
    .B(_00857_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05588_ (.A1(_00843_),
    .A2(_00849_),
    .A3(_00853_),
    .A4(_00857_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05589_ (.A1(_00842_),
    .A2(_00858_),
    .B(_00859_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05590_ (.A1(_00692_),
    .A2(_00702_),
    .A3(_00709_),
    .B(_00718_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05591_ (.A1(_00636_),
    .A2(_00762_),
    .A3(_00861_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05592_ (.A1(_00760_),
    .A2(_00776_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05593_ (.A1(_00760_),
    .A2(_00822_),
    .B1(_00863_),
    .B2(_00772_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05594_ (.A1(_00793_),
    .A2(_00862_),
    .A3(_00864_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05595_ (.A1(_00564_),
    .A2(_00855_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05596_ (.A1(_00787_),
    .A2(\as2650.instruction_args_latch[3] ),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05597_ (.A1(_00785_),
    .A2(_00866_),
    .B(_00867_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05598_ (.A1(_00865_),
    .A2(_00868_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05599_ (.I(_00794_),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05600_ (.A1(_00862_),
    .A2(_00864_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05601_ (.A1(_00870_),
    .A2(_00871_),
    .A3(_00868_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05602_ (.A1(_00860_),
    .A2(_00869_),
    .B(_00872_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05603_ (.A1(_00718_),
    .A2(_00740_),
    .A3(_00776_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05604_ (.A1(_00732_),
    .A2(_00874_),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05605_ (.A1(_00833_),
    .A2(_00875_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05606_ (.I(_00876_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05607_ (.A1(_00762_),
    .A2(_00765_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05608_ (.I(_00763_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05609_ (.A1(net262),
    .A2(_00764_),
    .B(_00879_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05610_ (.A1(_00879_),
    .A2(_00822_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05611_ (.A1(_00798_),
    .A2(_00878_),
    .A3(_00880_),
    .B(_00881_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05612_ (.I(_00882_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05613_ (.A1(_00561_),
    .A2(_00578_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05614_ (.A1(_00787_),
    .A2(_00814_),
    .A3(_00884_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05615_ (.A1(_00533_),
    .A2(\as2650.instruction_args_latch[5] ),
    .B(_00885_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05616_ (.A1(_00625_),
    .A2(_00877_),
    .A3(_00883_),
    .B(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05617_ (.A1(_00843_),
    .A2(_00876_),
    .A3(_00882_),
    .A4(_00886_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05618_ (.A1(_00574_),
    .A2(_00577_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05619_ (.A1(_00785_),
    .A2(_00578_),
    .A3(_00889_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05620_ (.A1(_00533_),
    .A2(\as2650.instruction_args_latch[4] ),
    .B(_00890_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05621_ (.A1(_00764_),
    .A2(_00761_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05622_ (.I(_00764_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05623_ (.A1(_00636_),
    .A2(_00893_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05624_ (.A1(_00637_),
    .A2(_00892_),
    .B(_00894_),
    .C(_00772_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05625_ (.A1(_00774_),
    .A2(_00776_),
    .B(_00741_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05626_ (.A1(_00896_),
    .A2(_00874_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05627_ (.A1(_00833_),
    .A2(_00897_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05628_ (.A1(_00625_),
    .A2(_00891_),
    .A3(_00895_),
    .A4(_00898_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05629_ (.I(_00895_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05630_ (.I(_00898_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05631_ (.A1(_00625_),
    .A2(_00900_),
    .A3(_00901_),
    .B(_00891_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _05632_ (.A1(_00887_),
    .A2(_00888_),
    .A3(_00899_),
    .A4(_00902_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05633_ (.A1(_00873_),
    .A2(_00903_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05634_ (.I(_00843_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _05635_ (.I(net238),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _05636_ (.A1(_00905_),
    .A2(_00906_),
    .A3(_00790_),
    .B1(_00813_),
    .B2(_00817_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05637_ (.A1(_00905_),
    .A2(_00906_),
    .B(_00790_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _05638_ (.A1(_00905_),
    .A2(_00877_),
    .A3(_00883_),
    .A4(_00886_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05639_ (.A1(_00905_),
    .A2(_00891_),
    .A3(_00900_),
    .A4(_00901_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05640_ (.A1(_00909_),
    .A2(_00910_),
    .B(_00887_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05641_ (.A1(_00791_),
    .A2(_00805_),
    .A3(net235),
    .A4(_00911_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _05642_ (.A1(_00820_),
    .A2(_00904_),
    .B1(_00907_),
    .B2(_00908_),
    .C(_00912_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05643_ (.A1(_00585_),
    .A2(_00587_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05644_ (.I(_00588_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05645_ (.A1(_00914_),
    .A2(_00915_),
    .B(_00599_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05646_ (.A1(_00534_),
    .A2(\as2650.instruction_args_latch[11] ),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05647_ (.A1(_00589_),
    .A2(_00916_),
    .B(_00917_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05648_ (.I(_00533_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05649_ (.A1(_00585_),
    .A2(_00587_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05650_ (.A1(_00919_),
    .A2(\as2650.instruction_args_latch[10] ),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05651_ (.A1(_00919_),
    .A2(_00914_),
    .A3(_00920_),
    .B(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05652_ (.A1(_00551_),
    .A2(_00579_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05653_ (.A1(_00923_),
    .A2(_00580_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05654_ (.A1(_00534_),
    .A2(\as2650.instruction_args_latch[8] ),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05655_ (.A1(_00534_),
    .A2(_00924_),
    .B(_00925_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05656_ (.A1(_00581_),
    .A2(_00584_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05657_ (.A1(_00919_),
    .A2(_00927_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05658_ (.A1(_00919_),
    .A2(\as2650.instruction_args_latch[9] ),
    .B1(_00585_),
    .B2(_00928_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05659_ (.I(_00929_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05660_ (.A1(_00918_),
    .A2(_00922_),
    .A3(_00926_),
    .A4(_00930_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05661_ (.I(_00931_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05662_ (.A1(_00589_),
    .A2(_00592_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05663_ (.A1(_00535_),
    .A2(_00933_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05664_ (.A1(_00535_),
    .A2(\as2650.instruction_args_latch[12] ),
    .B1(_00593_),
    .B2(_00934_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05665_ (.A1(net241),
    .A2(_00932_),
    .A3(_00935_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05666_ (.A1(_00629_),
    .A2(_00537_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05667_ (.I(_00599_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05668_ (.A1(\as2650.page_reg[1] ),
    .A2(_00528_),
    .B(_00938_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05669_ (.A1(\as2650.indirect_target[14] ),
    .A2(_00590_),
    .B1(_00594_),
    .B2(\as2650.page_reg[1] ),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05670_ (.A1(_00596_),
    .A2(_00940_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05671_ (.I(_00938_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05672_ (.A1(_00937_),
    .A2(_00939_),
    .B1(_00941_),
    .B2(_00942_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05673_ (.A1(_00601_),
    .A2(_00936_),
    .A3(_00943_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05674_ (.I(_00535_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05675_ (.A1(_00593_),
    .A2(_00595_),
    .A3(_00940_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05676_ (.A1(\as2650.indirect_target[15] ),
    .A2(_00590_),
    .B1(_00594_),
    .B2(\as2650.page_reg[2] ),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05677_ (.A1(_00946_),
    .A2(_00947_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05678_ (.I(\as2650.page_reg[2] ),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05679_ (.A1(_00949_),
    .A2(_00528_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05680_ (.A1(\as2650.instruction_args_latch[15] ),
    .A2(_00537_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05681_ (.A1(_00950_),
    .A2(_00951_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05682_ (.A1(_00945_),
    .A2(_00952_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05683_ (.A1(_00945_),
    .A2(_00948_),
    .B(_00953_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05684_ (.A1(_00944_),
    .A2(_00954_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05685_ (.A1(_00955_),
    .A2(\as2650.last_addr[15] ),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05686_ (.A1(_00540_),
    .A2(_00600_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _05687_ (.A1(_00957_),
    .A2(net241),
    .A3(_00932_),
    .A4(_00935_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05688_ (.A1(_00958_),
    .A2(_00943_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05689_ (.A1(\as2650.last_addr[14] ),
    .A2(_00959_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _05690_ (.A1(_00792_),
    .A2(_00806_),
    .A3(_00819_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05691_ (.A1(net243),
    .A2(_00903_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05692_ (.A1(_00792_),
    .A2(_00806_),
    .A3(_00819_),
    .A4(_00911_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05693_ (.A1(net250),
    .A2(_00908_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _05694_ (.A1(_00961_),
    .A2(_00962_),
    .B(_00963_),
    .C(_00964_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05695_ (.I(_00926_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05696_ (.A1(_00965_),
    .A2(_00966_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _05697_ (.A1(\as2650.last_addr[9] ),
    .A2(_00930_),
    .A3(_00967_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05698_ (.A1(net241),
    .A2(_00966_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05699_ (.A1(\as2650.last_addr[8] ),
    .A2(_00969_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05700_ (.A1(_00965_),
    .A2(_00931_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _05701_ (.A1(\as2650.last_addr[12] ),
    .A2(_00971_),
    .A3(_00935_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05702_ (.A1(_00968_),
    .A2(_00970_),
    .A3(_00972_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _05703_ (.A1(\as2650.last_addr[13] ),
    .A2(_00957_),
    .A3(_00936_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05704_ (.A1(_00965_),
    .A2(_00966_),
    .A3(_00930_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _05705_ (.A1(\as2650.last_addr[10] ),
    .A2(_00922_),
    .A3(_00975_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05706_ (.A1(_00974_),
    .A2(_00976_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05707_ (.A1(_00965_),
    .A2(_00922_),
    .A3(_00966_),
    .A4(_00930_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05708_ (.A1(_00918_),
    .A2(_00978_),
    .B(_00971_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _05709_ (.A1(\as2650.last_addr[11] ),
    .A2(_00979_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05710_ (.A1(_00960_),
    .A2(_00973_),
    .A3(_00977_),
    .A4(_00980_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05711_ (.A1(net237),
    .A2(_00888_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05712_ (.A1(_00899_),
    .A2(_00902_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05713_ (.A1(net244),
    .A2(_00983_),
    .B(_00910_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _05714_ (.A1(_00982_),
    .A2(_00984_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _05715_ (.A1(net384),
    .A2(_00869_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05716_ (.A1(_00849_),
    .A2(_00853_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05717_ (.A1(_00870_),
    .A2(_00987_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _05718_ (.A1(_00988_),
    .A2(_00857_),
    .A3(net257),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05719_ (.A1(_00870_),
    .A2(_00825_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _05720_ (.A1(_00990_),
    .A2(_00831_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05721_ (.A1(\as2650.last_addr[0] ),
    .A2(_00991_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05722_ (.A1(_00870_),
    .A2(_00840_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _05723_ (.A1(_00993_),
    .A2(_00838_),
    .A3(_00832_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05724_ (.A1(\as2650.last_addr[1] ),
    .A2(_00994_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05725_ (.A1(\as2650.last_addr[2] ),
    .A2(_00989_),
    .B(_00992_),
    .C(_00995_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _05726_ (.A1(\as2650.last_addr[3] ),
    .A2(_00986_),
    .B1(net258),
    .B2(\as2650.last_addr[2] ),
    .C(_00996_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05727_ (.A1(\as2650.last_addr[3] ),
    .A2(_00986_),
    .B(_00997_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _05728_ (.A1(net244),
    .A2(_00983_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05729_ (.A1(\as2650.last_addr[4] ),
    .A2(_00999_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05730_ (.A1(\as2650.last_addr[5] ),
    .A2(_00985_),
    .B(_00998_),
    .C(_01000_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05731_ (.A1(_00962_),
    .A2(_00911_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _05732_ (.A1(_00819_),
    .A2(_01002_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05733_ (.A1(\as2650.last_addr[6] ),
    .A2(_01003_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05734_ (.A1(\as2650.last_addr[5] ),
    .A2(_00985_),
    .B(_01001_),
    .C(_01004_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05735_ (.A1(_00792_),
    .A2(_00806_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05736_ (.A1(_00813_),
    .A2(_00817_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05737_ (.A1(_00813_),
    .A2(_00817_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05738_ (.A1(_01007_),
    .A2(_01002_),
    .B(_01008_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _05739_ (.A1(_01006_),
    .A2(_01009_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05740_ (.A1(\as2650.last_addr[7] ),
    .A2(_01010_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05741_ (.A1(_01011_),
    .A2(_01005_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _05742_ (.A1(\as2650.cycle[3] ),
    .A2(_00956_),
    .A3(_00981_),
    .A4(_01012_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05743_ (.A1(_01013_),
    .A2(_00530_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05744_ (.I(_01014_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05745_ (.I0(_00529_),
    .I1(\as2650.instruction_args_latch[15] ),
    .S(_01015_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05746_ (.I(_00613_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05747_ (.I(_01017_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05748_ (.I(_00602_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05749_ (.A1(_01018_),
    .A2(_01019_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05750_ (.A1(_00528_),
    .A2(_01016_),
    .B(_01020_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05751_ (.A1(_00521_),
    .A2(_01021_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05752_ (.I(net9),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05753_ (.A1(_01023_),
    .A2(_00516_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05754_ (.A1(\as2650.insin[3] ),
    .A2(_00516_),
    .B(_01024_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05755_ (.I(_01025_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05756_ (.I(_00603_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05757_ (.A1(_01026_),
    .A2(_01027_),
    .B(_00622_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05758_ (.I(_00526_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05759_ (.A1(_00524_),
    .A2(_01027_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05760_ (.A1(_01025_),
    .A2(_01030_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05761_ (.I(_01031_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05762_ (.A1(_01029_),
    .A2(_01032_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05763_ (.A1(_01028_),
    .A2(_01033_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05764_ (.I(_00956_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05765_ (.I(_00981_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05766_ (.A1(_01035_),
    .A2(_01036_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05767_ (.A1(_01011_),
    .A2(_01005_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05768_ (.A1(_01037_),
    .A2(_01038_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05769_ (.I(_01039_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05770_ (.I(_01040_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05771_ (.A1(_01022_),
    .A2(_01034_),
    .B(_01041_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05772_ (.I(_01026_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05773_ (.I(_01012_),
    .Z(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05774_ (.A1(_00565_),
    .A2(_01035_),
    .A3(_01036_),
    .A4(_01044_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05775_ (.I(_01045_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05776_ (.A1(_00528_),
    .A2(_01016_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05777_ (.I(_01047_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05778_ (.A1(_01043_),
    .A2(_01046_),
    .A3(_01048_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05779_ (.I(_01049_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05780_ (.A1(_00512_),
    .A2(_01042_),
    .B(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05781_ (.I(_00530_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05782_ (.I(_01052_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05783_ (.I(_01053_),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05784_ (.A1(_01054_),
    .A2(_01039_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05785_ (.I(_00517_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05786_ (.I(_01056_),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05787_ (.I(_01057_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05788_ (.I(_01058_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05789_ (.I(_00770_),
    .Z(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05790_ (.I(net4),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05791_ (.A1(_01061_),
    .A2(_00517_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05792_ (.A1(\as2650.insin[7] ),
    .A2(_01056_),
    .B(_01062_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05793_ (.I(net3),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05794_ (.I(_01064_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05795_ (.A1(_01065_),
    .A2(_00517_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05796_ (.A1(\as2650.insin[6] ),
    .A2(_01056_),
    .B(_01066_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05797_ (.A1(_01063_),
    .A2(_01067_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05798_ (.A1(_00613_),
    .A2(_01068_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05799_ (.I(_01069_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05800_ (.I(_00608_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05801_ (.A1(_01071_),
    .A2(_01069_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05802_ (.I(_01072_),
    .Z(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05803_ (.A1(_00800_),
    .A2(_00801_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05804_ (.A1(_00613_),
    .A2(_01068_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05805_ (.A1(_01071_),
    .A2(_01075_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05806_ (.A1(_00751_),
    .A2(_00768_),
    .B(_01076_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _05807_ (.A1(_01060_),
    .A2(_01070_),
    .B1(_01073_),
    .B2(_01074_),
    .C(_01077_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05808_ (.I(_00773_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05809_ (.I(net2),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05810_ (.A1(_01080_),
    .A2(_01056_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05811_ (.A1(\as2650.insin[5] ),
    .A2(_01057_),
    .B(_01081_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05812_ (.I(_01082_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05813_ (.A1(_01083_),
    .A2(_01070_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05814_ (.A1(_00807_),
    .A2(_00808_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05815_ (.A1(_01079_),
    .A2(_01070_),
    .B1(_01073_),
    .B2(net249),
    .C1(_01084_),
    .C2(_01085_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05816_ (.I(_00732_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05817_ (.I(_01075_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05818_ (.A1(_01083_),
    .A2(_01075_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05819_ (.A1(_00878_),
    .A2(_00880_),
    .A3(_01076_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05820_ (.A1(_01087_),
    .A2(_01088_),
    .B1(_01089_),
    .B2(net382),
    .C(_01090_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05821_ (.A1(_00762_),
    .A2(_00861_),
    .A3(_01084_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05822_ (.I(_00760_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05823_ (.A1(_01093_),
    .A2(_01070_),
    .B1(_01073_),
    .B2(_00863_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05824_ (.A1(_01092_),
    .A2(_01094_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05825_ (.I(_00741_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _05826_ (.A1(_01096_),
    .A2(_01088_),
    .B1(_01089_),
    .B2(net261),
    .C1(_01076_),
    .C2(net253),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05827_ (.A1(_00845_),
    .A2(_00846_),
    .B(_00848_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05828_ (.A1(_01098_),
    .A2(_01084_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05829_ (.A1(_00846_),
    .A2(_01088_),
    .B1(_01089_),
    .B2(_00851_),
    .C(_01099_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05830_ (.I(_00844_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05831_ (.A1(_01101_),
    .A2(_01088_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05832_ (.A1(_00845_),
    .A2(_00850_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05833_ (.A1(_00844_),
    .A2(_01076_),
    .B(_01072_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05834_ (.A1(_01103_),
    .A2(_01104_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05835_ (.A1(_01097_),
    .A2(_01100_),
    .A3(_01102_),
    .A4(_01105_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05836_ (.A1(_01091_),
    .A2(_01095_),
    .A3(_01106_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05837_ (.I(_01067_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05838_ (.A1(_01017_),
    .A2(_01108_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05839_ (.A1(_01078_),
    .A2(_01086_),
    .A3(_01107_),
    .B(_01109_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05840_ (.I(_01019_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05841_ (.I(_00524_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05842_ (.I(_00610_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05843_ (.I(_01113_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05844_ (.A1(_01017_),
    .A2(_01108_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05845_ (.A1(_01114_),
    .A2(_01115_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05846_ (.A1(_01112_),
    .A2(_00645_),
    .A3(_01116_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05847_ (.I(_00610_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05848_ (.A1(_01118_),
    .A2(_01109_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05849_ (.I(_01119_),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05850_ (.I(_00641_),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05851_ (.A1(\as2650.debug_psl[6] ),
    .A2(_01121_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05852_ (.A1(\as2650.debug_psl[6] ),
    .A2(_01121_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05853_ (.A1(\as2650.debug_psl[7] ),
    .A2(_00639_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05854_ (.A1(_01122_),
    .A2(_01123_),
    .B(_01124_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05855_ (.I(_01125_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05856_ (.A1(_00645_),
    .A2(_01126_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05857_ (.A1(_01116_),
    .A2(_01125_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _05858_ (.A1(_01111_),
    .A2(_01117_),
    .B1(_01120_),
    .B2(_01127_),
    .C(_01128_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _05859_ (.A1(_00614_),
    .A2(_01110_),
    .A3(_01129_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05860_ (.I(_01130_),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05861_ (.I(_01131_),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05862_ (.I(_01132_),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05863_ (.I(_00645_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05864_ (.I(_01018_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05865_ (.A1(_01112_),
    .A2(_01019_),
    .A3(_00520_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05866_ (.A1(_01135_),
    .A2(_01136_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05867_ (.I(_01071_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05868_ (.A1(_01063_),
    .A2(_00611_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05869_ (.A1(_01138_),
    .A2(_01139_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05870_ (.I(_01140_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05871_ (.A1(_01134_),
    .A2(_01137_),
    .A3(_01141_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05872_ (.A1(_01082_),
    .A2(_01139_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05873_ (.I(_01143_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05874_ (.A1(_01137_),
    .A2(_01144_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05875_ (.I(_00606_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05876_ (.I(_01146_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05877_ (.I(_00611_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05878_ (.A1(_00610_),
    .A2(_01148_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05879_ (.A1(_00609_),
    .A2(_01149_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05880_ (.A1(_01120_),
    .A2(_01150_),
    .B(_01136_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05881_ (.A1(_01025_),
    .A2(_00520_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05882_ (.I(_01152_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05883_ (.I(_01153_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05884_ (.I(_01154_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05885_ (.I(_01155_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05886_ (.A1(_01147_),
    .A2(_00604_),
    .A3(_01151_),
    .A4(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05887_ (.A1(_01142_),
    .A2(_01145_),
    .A3(_01157_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05888_ (.A1(_01032_),
    .A2(_01158_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05889_ (.I(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05890_ (.I(_01160_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05891_ (.A1(_01059_),
    .A2(_01133_),
    .A3(_01161_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05892_ (.A1(_00510_),
    .A2(_01051_),
    .B1(_01055_),
    .B2(_01162_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05893_ (.I(_00509_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05894_ (.I(_01041_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05895_ (.A1(_01043_),
    .A2(_01048_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05896_ (.I(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _05897_ (.A1(\as2650.last_addr[15] ),
    .A2(_00955_),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05898_ (.A1(_00960_),
    .A2(_00973_),
    .A3(_00977_),
    .A4(_00980_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05899_ (.A1(_00566_),
    .A2(_01167_),
    .A3(_01168_),
    .A4(_01038_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05900_ (.A1(_00530_),
    .A2(_01169_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05901_ (.I(_01170_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05902_ (.I(_01171_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05903_ (.I(_01172_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _05904_ (.A1(_00942_),
    .A2(_01163_),
    .A3(_01164_),
    .B1(_01166_),
    .B2(_01173_),
    .B3(_00614_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05905_ (.I(_01015_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05906_ (.I(_01028_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05907_ (.I(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05908_ (.I(_01176_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05909_ (.I(_00565_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05910_ (.I(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05911_ (.I(_01053_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05912_ (.I(_01180_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05913_ (.I(_01181_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05914_ (.I(_01182_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05915_ (.I(_01183_),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05916_ (.A1(_01035_),
    .A2(_01036_),
    .A3(_01044_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05917_ (.I(_01185_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05918_ (.I(_01186_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05919_ (.A1(_01179_),
    .A2(_01184_),
    .A3(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05920_ (.A1(_01174_),
    .A2(_01177_),
    .A3(_01033_),
    .B(_01188_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05921_ (.I(_01021_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05922_ (.A1(_01022_),
    .A2(_01033_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05923_ (.A1(_01176_),
    .A2(_01190_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05924_ (.A1(_01178_),
    .A2(_01189_),
    .B1(_01191_),
    .B2(_00511_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05925_ (.I(_01192_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05926_ (.A1(_01032_),
    .A2(_01158_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05927_ (.I(_01194_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05928_ (.I(_01195_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05929_ (.I(_01108_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05930_ (.A1(_01113_),
    .A2(_01197_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05931_ (.I(_00654_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05932_ (.I(_01199_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05933_ (.I(_01200_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05934_ (.I(_01201_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05935_ (.A1(_01026_),
    .A2(_01030_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05936_ (.A1(_00609_),
    .A2(_01202_),
    .A3(_01203_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05937_ (.A1(_01198_),
    .A2(_01204_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05938_ (.I(_01205_),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05939_ (.I(_01135_),
    .Z(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05940_ (.I(_01138_),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05941_ (.A1(_00524_),
    .A2(_01019_),
    .A3(_01027_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05942_ (.I(_01209_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _05943_ (.A1(_01207_),
    .A2(_01208_),
    .A3(_01210_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05944_ (.A1(_01196_),
    .A2(_01206_),
    .A3(_01211_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05945_ (.I(_01057_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05946_ (.I(_01213_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05947_ (.A1(_01133_),
    .A2(_01212_),
    .B(_01214_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05948_ (.A1(_01193_),
    .A2(_01215_),
    .B(_01164_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05949_ (.A1(_00945_),
    .A2(_01040_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05950_ (.A1(_01182_),
    .A2(_01217_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05951_ (.I(_01218_),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05952_ (.A1(_01059_),
    .A2(_01187_),
    .B(_01219_),
    .C(\as2650.cycle[4] ),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05953_ (.A1(_01216_),
    .A2(_01220_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05954_ (.A1(_00647_),
    .A2(\as2650.regs[0][0] ),
    .Z(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05955_ (.A1(_00727_),
    .A2(\as2650.regs[4][0] ),
    .B(_01221_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05956_ (.I(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05957_ (.I(_01223_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05958_ (.I(_01224_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05959_ (.I(_01225_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05960_ (.I(_01226_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05961_ (.I(_01227_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05962_ (.I(_01228_),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05963_ (.A1(_00648_),
    .A2(\as2650.regs[0][1] ),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05964_ (.A1(_00671_),
    .A2(\as2650.regs[4][1] ),
    .B(_01229_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05965_ (.I(_01230_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05966_ (.I(_01231_),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05967_ (.I(_01232_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05968_ (.I(_01233_),
    .Z(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05969_ (.I(_01234_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05970_ (.I(_01235_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05971_ (.I(_01236_),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05972_ (.A1(_00648_),
    .A2(\as2650.regs[0][2] ),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05973_ (.A1(_00671_),
    .A2(\as2650.regs[4][2] ),
    .B(_01237_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05974_ (.I(_01238_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05975_ (.I(_01239_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05976_ (.I(_01240_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05977_ (.I(_01241_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05978_ (.I(_01242_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05979_ (.I(_01243_),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05980_ (.I(_00736_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05981_ (.A1(_00710_),
    .A2(\as2650.regs[0][3] ),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05982_ (.A1(_01244_),
    .A2(\as2650.regs[4][3] ),
    .B(_01245_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05983_ (.I(_01246_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05984_ (.I(_01247_),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05985_ (.I(_01248_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05986_ (.I(_01249_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05987_ (.I(_01250_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05988_ (.I(_01251_),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05989_ (.A1(_00647_),
    .A2(\as2650.regs[0][4] ),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05990_ (.A1(_00736_),
    .A2(\as2650.regs[4][4] ),
    .B(_01252_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05991_ (.I(_01253_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05992_ (.I(_01254_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05993_ (.I(_01255_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05994_ (.I(_01256_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05995_ (.I(_01257_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05996_ (.I(_01258_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05997_ (.I(_01259_),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05998_ (.A1(_00649_),
    .A2(\as2650.regs[0][5] ),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05999_ (.A1(_00746_),
    .A2(\as2650.regs[4][5] ),
    .B(_01260_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06000_ (.I(_01261_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06001_ (.I(_01262_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06002_ (.I(_01263_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06003_ (.I(_01264_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06004_ (.I(_01265_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06005_ (.I(_01266_),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06006_ (.A1(_00649_),
    .A2(\as2650.regs[0][6] ),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06007_ (.A1(_00746_),
    .A2(\as2650.regs[4][6] ),
    .B(_01267_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06008_ (.I(_01268_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06009_ (.I(_01269_),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06010_ (.I(_01270_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06011_ (.I(_01271_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06012_ (.I(_01272_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06013_ (.I(_01273_),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06014_ (.A1(_00672_),
    .A2(\as2650.regs[4][7] ),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06015_ (.A1(_00650_),
    .A2(\as2650.regs[0][7] ),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06016_ (.A1(_01274_),
    .A2(_01275_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06017_ (.I(_01276_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06018_ (.I(_01277_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06019_ (.I(_01278_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06020_ (.I(_01279_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06021_ (.I(_01280_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06022_ (.I(_01281_),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06023_ (.A1(\as2650.cycle[4] ),
    .A2(\as2650.cycle[1] ),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06024_ (.A1(_01018_),
    .A2(_01208_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06025_ (.A1(_01203_),
    .A2(_01283_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06026_ (.A1(\as2650.cycle[1] ),
    .A2(_01114_),
    .A3(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06027_ (.A1(_00622_),
    .A2(_00511_),
    .B(_00945_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06028_ (.A1(_00609_),
    .A2(_01149_),
    .A3(_01204_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06029_ (.A1(_01146_),
    .A2(_01111_),
    .B(_01287_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06030_ (.I(_01288_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06031_ (.A1(_01286_),
    .A2(_01289_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06032_ (.A1(_01186_),
    .A2(_01282_),
    .B1(_01285_),
    .B2(_01290_),
    .C(_00508_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06033_ (.A1(_00546_),
    .A2(_00567_),
    .B(\as2650.cycle[4] ),
    .C(\as2650.cycle[1] ),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06034_ (.A1(_01035_),
    .A2(_01036_),
    .A3(_01038_),
    .A4(_01292_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06035_ (.I(_01293_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06036_ (.I(_01294_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06037_ (.A1(_01037_),
    .A2(_01292_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06038_ (.I(_01296_),
    .Z(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06039_ (.I(_01063_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06040_ (.A1(_01298_),
    .A2(_01211_),
    .A3(_01282_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06041_ (.I(_01299_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06042_ (.A1(_01295_),
    .A2(_01297_),
    .A3(_01300_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06043_ (.I(_01182_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06044_ (.I(_01302_),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06045_ (.I(_01303_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06046_ (.A1(_01291_),
    .A2(_01301_),
    .B(_01304_),
    .ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06047_ (.I(_01185_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06048_ (.A1(_00546_),
    .A2(_00567_),
    .B(_01305_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06049_ (.A1(_01114_),
    .A2(_01211_),
    .A3(_01282_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06050_ (.I(_01302_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06051_ (.A1(_01306_),
    .A2(_01307_),
    .B(_01308_),
    .C(_01290_),
    .ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06052_ (.I(_01296_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06053_ (.I(_01309_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06054_ (.A1(clknet_leaf_27_wb_clk_i),
    .A2(_01184_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06055_ (.A1(_01310_),
    .A2(clknet_1_0__leaf__01311_),
    .ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06056_ (.I(_01293_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06057_ (.I(_01312_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06058_ (.A1(_01313_),
    .A2(clknet_1_1__leaf__01311_),
    .ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06059_ (.A1(\web_behavior[1] ),
    .A2(clknet_leaf_107_wb_clk_i),
    .B(\web_behavior[0] ),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06060_ (.A1(\web_behavior[1] ),
    .A2(clknet_leaf_108_wb_clk_i),
    .B(\web_behavior[0] ),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06061__1 (.I(_01315_),
    .ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06062_ (.A1(_01314_),
    .A2(net231),
    .B(_01291_),
    .ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06063_ (.I(wb_debug_carry),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06064_ (.I(\as2650.debug_psl[0] ),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06065_ (.I(\as2650.debug_psl[6] ),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06066_ (.I(_01319_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06067_ (.I(_01148_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06068_ (.A1(wb_debug_cc),
    .A2(_01282_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06069_ (.A1(wb_debug_cc),
    .A2(_01320_),
    .B1(_01321_),
    .B2(_01322_),
    .C(_01317_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06070_ (.A1(_01317_),
    .A2(_01318_),
    .B(_01323_),
    .ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06071_ (.I(\as2650.debug_psl[5] ),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06072_ (.I(_01324_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06073_ (.I(\as2650.debug_psl[7] ),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06074_ (.I(_01326_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06075_ (.I(_01197_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06076_ (.A1(wb_debug_cc),
    .A2(_01327_),
    .B1(_01328_),
    .B2(_01322_),
    .C(wb_debug_carry),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06077_ (.A1(_01317_),
    .A2(_01325_),
    .B(_01329_),
    .ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06078_ (.I0(\as2650.regs[1][5] ),
    .I1(\as2650.regs[5][5] ),
    .S(_00727_),
    .Z(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06079_ (.I(_01330_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06080_ (.I(_01331_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06081_ (.I(_01332_),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06082_ (.I0(\as2650.regs[1][4] ),
    .I1(\as2650.regs[5][4] ),
    .S(_00671_),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06083_ (.I(_01333_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06084_ (.I(_01334_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06085_ (.I(_01335_),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06086_ (.I0(\as2650.regs[1][3] ),
    .I1(\as2650.regs[5][3] ),
    .S(_01244_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06087_ (.I(_01336_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06088_ (.I(_01337_),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06089_ (.I(_01338_),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06090_ (.I0(\as2650.regs[1][2] ),
    .I1(\as2650.regs[5][2] ),
    .S(_01244_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06091_ (.I(_01339_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06092_ (.I(_01340_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06093_ (.I(_01341_),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06094_ (.I0(\as2650.regs[1][6] ),
    .I1(\as2650.regs[5][6] ),
    .S(_01244_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06095_ (.I(_01342_),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06096_ (.I(_01343_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06097_ (.I(_01344_),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06098_ (.I0(\as2650.regs[1][1] ),
    .I1(\as2650.regs[5][1] ),
    .S(_00672_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06099_ (.I(_01345_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06100_ (.I(_01346_),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06101_ (.I(_01347_),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06102_ (.I(_01348_),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06103_ (.I(_00672_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06104_ (.I0(\as2650.regs[1][0] ),
    .I1(\as2650.regs[5][0] ),
    .S(_01349_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06105_ (.I(_01350_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06106_ (.I(_01351_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06107_ (.I(_01352_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06108_ (.I(_01353_),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06109_ (.I0(\as2650.regs[1][7] ),
    .I1(\as2650.regs[5][7] ),
    .S(_00677_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06110_ (.I(_01354_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06111_ (.I(_01355_),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06112_ (.I(_01349_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06113_ (.I(_01356_),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06114_ (.I(_01357_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06115_ (.I(_01358_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06116_ (.I(_01359_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06117_ (.I(_01360_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06118_ (.I(_01361_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06119_ (.I0(\as2650.regs[2][0] ),
    .I1(\as2650.regs[6][0] ),
    .S(_01362_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06120_ (.I(_01363_),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06121_ (.I0(\as2650.regs[2][1] ),
    .I1(\as2650.regs[6][1] ),
    .S(_01362_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06122_ (.I(_01364_),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06123_ (.I0(\as2650.regs[2][2] ),
    .I1(\as2650.regs[6][2] ),
    .S(_01362_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06124_ (.I(_01365_),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06125_ (.I0(\as2650.regs[2][3] ),
    .I1(\as2650.regs[6][3] ),
    .S(_01362_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06126_ (.I(_01366_),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06127_ (.I(_01360_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06128_ (.I(_01367_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06129_ (.I(\as2650.regs[2][4] ),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06130_ (.A1(_01368_),
    .A2(\as2650.regs[6][4] ),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06131_ (.A1(_01368_),
    .A2(_01369_),
    .B(_01370_),
    .ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06132_ (.I(\as2650.regs[2][5] ),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06133_ (.A1(_01368_),
    .A2(\as2650.regs[6][5] ),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06134_ (.A1(_01368_),
    .A2(_01371_),
    .B(_01372_),
    .ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06135_ (.I0(\as2650.regs[2][6] ),
    .I1(\as2650.regs[6][6] ),
    .S(_01367_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06136_ (.I(_01373_),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06137_ (.I0(\as2650.regs[2][7] ),
    .I1(\as2650.regs[6][7] ),
    .S(_01367_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06138_ (.I(_01374_),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06139_ (.I0(\as2650.regs[3][0] ),
    .I1(\as2650.regs[7][0] ),
    .S(_01349_),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06140_ (.I(_01375_),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06141_ (.I0(\as2650.regs[3][1] ),
    .I1(\as2650.regs[7][1] ),
    .S(_01356_),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06142_ (.I(_01376_),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06143_ (.I0(\as2650.regs[3][2] ),
    .I1(\as2650.regs[7][2] ),
    .S(_01356_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06144_ (.I(_01377_),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06145_ (.I0(\as2650.regs[3][3] ),
    .I1(\as2650.regs[7][3] ),
    .S(_01356_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06146_ (.I(_01378_),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06147_ (.I0(\as2650.regs[3][4] ),
    .I1(\as2650.regs[7][4] ),
    .S(_01357_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06148_ (.I(_01379_),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06149_ (.I0(\as2650.regs[3][5] ),
    .I1(\as2650.regs[7][5] ),
    .S(_01357_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06150_ (.I(_01380_),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06151_ (.I0(\as2650.regs[3][6] ),
    .I1(\as2650.regs[7][6] ),
    .S(_01357_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06152_ (.I(_01381_),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06153_ (.I0(\as2650.regs[3][7] ),
    .I1(\as2650.regs[7][7] ),
    .S(_01358_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06154_ (.I(_01382_),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06155_ (.I(_01082_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06156_ (.I(_01383_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06157_ (.A1(_00602_),
    .A2(_00603_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06158_ (.I(_01385_),
    .Z(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06159_ (.I(_01386_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06160_ (.I(_01387_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06161_ (.I(_01388_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06162_ (.I(_01389_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06163_ (.I(_01390_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06164_ (.A1(_01384_),
    .A2(_01120_),
    .A3(_01391_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06165_ (.I(_01392_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06166_ (.A1(_01147_),
    .A2(_01134_),
    .A3(_01393_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06167_ (.A1(_01058_),
    .A2(_01040_),
    .A3(_01206_),
    .A4(_01394_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06168_ (.I(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06169_ (.A1(\as2650.chirp_ptr[1] ),
    .A2(\as2650.chirp_ptr[0] ),
    .A3(_01396_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06170_ (.A1(\as2650.chirp_ptr[2] ),
    .A2(_01397_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06171_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01396_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06172_ (.A1(_01181_),
    .A2(_01399_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06173_ (.I(_01400_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06174_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01396_),
    .B(\as2650.chirp_ptr[1] ),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06175_ (.A1(_01181_),
    .A2(_01397_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06176_ (.A1(_01401_),
    .A2(_01402_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06177_ (.I(_01403_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06178_ (.A1(_00210_),
    .A2(_00211_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06179_ (.A1(_01399_),
    .A2(_00211_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06180_ (.A1(_01404_),
    .A2(_01405_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06181_ (.A1(_00507_),
    .A2(_01398_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06182_ (.I(_01407_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06183_ (.A1(_01398_),
    .A2(_00210_),
    .B1(_01406_),
    .B2(_00212_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06184_ (.I(_01405_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06185_ (.I(_00212_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06186_ (.A1(_01409_),
    .A2(_01404_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06187_ (.A1(_01408_),
    .A2(_01410_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06188_ (.I(_01398_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06189_ (.A1(_01411_),
    .A2(_00211_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06190_ (.A1(_00212_),
    .A2(_01406_),
    .B(_01412_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06191_ (.A1(_01409_),
    .A2(_01404_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06192_ (.A1(_01409_),
    .A2(_01408_),
    .B(_01413_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06193_ (.A1(_01410_),
    .A2(_01412_),
    .Z(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06194_ (.I(_01414_),
    .Z(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06195_ (.I(_01299_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06196_ (.I(_01415_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06197_ (.A1(_00969_),
    .A2(_01297_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06198_ (.A1(_01037_),
    .A2(_01292_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06199_ (.I(_01418_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06200_ (.I(_01419_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06201_ (.A1(_01199_),
    .A2(_01227_),
    .B(_00938_),
    .C(_00619_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06202_ (.A1(_01199_),
    .A2(net255),
    .A3(_00824_),
    .B(_01421_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06203_ (.A1(_00621_),
    .A2(_00844_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06204_ (.A1(_01422_),
    .A2(_01423_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06205_ (.I(_01424_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06206_ (.A1(_01420_),
    .A2(_01425_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06207_ (.I(_01312_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06208_ (.A1(_01417_),
    .A2(_01426_),
    .B(_01427_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06209_ (.I(_01312_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06210_ (.I(_01429_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06211_ (.I(_01299_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06212_ (.A1(_00991_),
    .A2(_01430_),
    .B(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06213_ (.A1(_01101_),
    .A2(_01416_),
    .B1(_01428_),
    .B2(_01432_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06214_ (.I(_00755_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06215_ (.I(_01433_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06216_ (.I(_01415_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06217_ (.I(_01418_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06218_ (.I(_00670_),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06219_ (.I(_00692_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06220_ (.A1(_01438_),
    .A2(_00847_),
    .A3(_00834_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06221_ (.A1(_00938_),
    .A2(_00619_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06222_ (.I(_01199_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06223_ (.I(_01230_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06224_ (.A1(_01441_),
    .A2(_01442_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06225_ (.A1(_01440_),
    .A2(_01443_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06226_ (.A1(_01437_),
    .A2(_01439_),
    .B(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06227_ (.I(_01440_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06228_ (.A1(_01446_),
    .A2(_00755_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06229_ (.A1(_01445_),
    .A2(_01447_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06230_ (.I(_01448_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06231_ (.A1(_00929_),
    .A2(_00967_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06232_ (.A1(_00975_),
    .A2(_01450_),
    .A3(_01419_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06233_ (.A1(_01436_),
    .A2(_01449_),
    .B(_01451_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06234_ (.I(_01312_),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06235_ (.A1(_00994_),
    .A2(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06236_ (.A1(_01427_),
    .A2(_01452_),
    .B(_01454_),
    .C(_01415_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06237_ (.A1(_01434_),
    .A2(_01435_),
    .B(_01455_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06238_ (.I(_00759_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06239_ (.I(_01456_),
    .Z(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06240_ (.A1(_00922_),
    .A2(_00975_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06241_ (.A1(_01458_),
    .A2(_01297_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06242_ (.I(_00621_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06243_ (.A1(_01441_),
    .A2(_01243_),
    .B(_01460_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06244_ (.A1(_01441_),
    .A2(_00849_),
    .A3(_00853_),
    .B(_01461_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06245_ (.A1(_01460_),
    .A2(_01456_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06246_ (.A1(_01462_),
    .A2(_01463_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06247_ (.I(_01464_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06248_ (.A1(_01420_),
    .A2(_01465_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06249_ (.A1(_01459_),
    .A2(_01466_),
    .B(_01427_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06250_ (.A1(_00989_),
    .A2(_01453_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06251_ (.A1(_01431_),
    .A2(_01468_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06252_ (.A1(_01457_),
    .A2(_01416_),
    .B1(_01467_),
    .B2(_01469_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06253_ (.I(_01093_),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06254_ (.I(_01446_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06255_ (.I(_00774_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06256_ (.A1(_00670_),
    .A2(_00862_),
    .A3(_00864_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06257_ (.A1(_01441_),
    .A2(_01251_),
    .B(_01460_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06258_ (.A1(_01473_),
    .A2(_01474_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06259_ (.A1(_01471_),
    .A2(_01472_),
    .B(_01475_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06260_ (.A1(_00979_),
    .A2(_01296_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06261_ (.A1(_01436_),
    .A2(_01476_),
    .B(_01477_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06262_ (.A1(_00986_),
    .A2(_01294_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06263_ (.A1(_01453_),
    .A2(_01478_),
    .B(_01479_),
    .C(_01415_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06264_ (.A1(_01470_),
    .A2(_01435_),
    .B(_01480_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06265_ (.A1(_01200_),
    .A2(_00900_),
    .A3(_00901_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06266_ (.I(_01253_),
    .Z(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06267_ (.A1(_01437_),
    .A2(_01482_),
    .B(_01446_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06268_ (.A1(_01446_),
    .A2(_01096_),
    .B1(_01481_),
    .B2(_01483_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06269_ (.I(_01484_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06270_ (.A1(_00971_),
    .A2(_00935_),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06271_ (.A1(_01486_),
    .A2(_01419_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06272_ (.A1(_01436_),
    .A2(_01485_),
    .B(_01487_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06273_ (.A1(_00999_),
    .A2(_01429_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06274_ (.A1(_01300_),
    .A2(_01489_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06275_ (.A1(_01295_),
    .A2(_01488_),
    .B(_01490_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06276_ (.A1(_00893_),
    .A2(_01435_),
    .B(_01491_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06277_ (.I(_00879_),
    .Z(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06278_ (.I(_00621_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06279_ (.A1(_01200_),
    .A2(_00877_),
    .A3(_00883_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06280_ (.A1(_01201_),
    .A2(_01266_),
    .B(_01493_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06281_ (.A1(_01493_),
    .A2(_00879_),
    .B1(_01494_),
    .B2(_01495_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06282_ (.I(_01496_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06283_ (.A1(_00601_),
    .A2(_00936_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06284_ (.A1(_01498_),
    .A2(_01419_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06285_ (.A1(_01436_),
    .A2(_01497_),
    .B(_01499_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06286_ (.A1(_00985_),
    .A2(_01294_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06287_ (.A1(_01453_),
    .A2(_01500_),
    .B(_01501_),
    .C(_01299_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06288_ (.A1(_01492_),
    .A2(_01435_),
    .B(_01502_),
    .ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06289_ (.I(_01079_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06290_ (.I(_01503_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06291_ (.I(_01504_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06292_ (.A1(_00959_),
    .A2(_01309_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06293_ (.I(_01493_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06294_ (.I(_00811_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06295_ (.I0(_00810_),
    .I1(_01508_),
    .S(_00632_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06296_ (.A1(_01437_),
    .A2(_01509_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06297_ (.A1(_01201_),
    .A2(_01271_),
    .B(_01507_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06298_ (.A1(_01507_),
    .A2(_00773_),
    .B1(_01510_),
    .B2(_01511_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06299_ (.I(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06300_ (.A1(_01420_),
    .A2(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06301_ (.A1(_01506_),
    .A2(_01514_),
    .B(_01427_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06302_ (.A1(_01003_),
    .A2(_01429_),
    .B(_01431_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06303_ (.A1(_01505_),
    .A2(_01416_),
    .B1(_01515_),
    .B2(_01516_),
    .ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06304_ (.I(_01060_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06305_ (.A1(_01201_),
    .A2(_01279_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06306_ (.A1(_01202_),
    .A2(_00906_),
    .B(_01518_),
    .C(_01471_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06307_ (.A1(_01471_),
    .A2(_00795_),
    .B(_01519_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06308_ (.I(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06309_ (.A1(_00955_),
    .A2(_01309_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06310_ (.A1(_01420_),
    .A2(_01521_),
    .B(_01522_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06311_ (.A1(_01295_),
    .A2(_01523_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06312_ (.A1(_01010_),
    .A2(_01429_),
    .B(_01431_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06313_ (.A1(_01517_),
    .A2(_01416_),
    .B1(_01524_),
    .B2(_01525_),
    .ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06314_ (.A1(\as2650.cycle[1] ),
    .A2(_01308_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06315_ (.I(_01526_),
    .Z(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06316_ (.I(_01206_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06317_ (.A1(_01214_),
    .A2(_01055_),
    .A3(_01527_),
    .A4(_01211_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06318_ (.I(_01528_),
    .Z(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06319_ (.I(_00509_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06320_ (.A1(\as2650.cycle[3] ),
    .A2(_00956_),
    .A3(net233),
    .A4(_01044_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06321_ (.I(_01530_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06322_ (.I(_01531_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06323_ (.A1(_01532_),
    .A2(_01034_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06324_ (.I(_01533_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06325_ (.A1(_01111_),
    .A2(_00521_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06326_ (.A1(_01207_),
    .A2(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06327_ (.A1(_01047_),
    .A2(_01536_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06328_ (.I(_01537_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06329_ (.I(_01013_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06330_ (.I(_01539_),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06331_ (.I(_01540_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06332_ (.A1(_01058_),
    .A2(_01541_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06333_ (.I(_01542_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06334_ (.A1(_01534_),
    .A2(_01538_),
    .B1(_01543_),
    .B2(_00622_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06335_ (.A1(_01529_),
    .A2(_01544_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06336_ (.I(net11),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06337_ (.I(wb_feedback_delay),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06338_ (.A1(_01545_),
    .A2(_01546_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06339_ (.I(net13),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06340_ (.I(_01547_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06341_ (.I(_01548_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06342_ (.I(\wb_counter[0] ),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06343_ (.A1(net12),
    .A2(_01547_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06344_ (.I(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06345_ (.I(_01552_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06346_ (.I(\as2650.debug_psl[0] ),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06347_ (.I(_01554_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06348_ (.I(_01555_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06349_ (.A1(net47),
    .A2(net14),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06350_ (.A1(wb_feedback_delay),
    .A2(_01557_),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06351_ (.I(_01558_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06352_ (.I(_01559_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06353_ (.I(_01560_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06354_ (.A1(_01549_),
    .A2(_01550_),
    .B1(_01553_),
    .B2(_01556_),
    .C(_01561_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06355_ (.A1(net47),
    .A2(net14),
    .A3(_01546_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06356_ (.I(_01563_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06357_ (.I(_01564_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06358_ (.A1(net107),
    .A2(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06359_ (.I(_01545_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06360_ (.A1(_01562_),
    .A2(_01566_),
    .B(_01567_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06361_ (.I(\as2650.debug_psl[1] ),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06362_ (.I(_01568_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06363_ (.I(_01552_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06364_ (.A1(_01549_),
    .A2(\wb_counter[1] ),
    .B1(_01569_),
    .B2(_01570_),
    .C(_01561_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06365_ (.A1(net118),
    .A2(_01565_),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06366_ (.A1(_01571_),
    .A2(_01572_),
    .B(_01567_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06367_ (.I(\as2650.debug_psl[2] ),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06368_ (.I(_01573_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06369_ (.A1(_01549_),
    .A2(\wb_counter[2] ),
    .B1(_01574_),
    .B2(_01570_),
    .C(_01561_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06370_ (.A1(net129),
    .A2(_01565_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06371_ (.A1(_01575_),
    .A2(_01576_),
    .B(_01567_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06372_ (.I(\as2650.debug_psl[3] ),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06373_ (.I(_01577_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06374_ (.I(_01578_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06375_ (.A1(_01549_),
    .A2(\wb_counter[3] ),
    .B1(_01579_),
    .B2(_01570_),
    .C(_01561_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06376_ (.A1(net132),
    .A2(_01565_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06377_ (.A1(_01580_),
    .A2(_01581_),
    .B(_01567_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06378_ (.I(_01548_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06379_ (.I(\wb_counter[4] ),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06380_ (.I(_01552_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06381_ (.I(_01560_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06382_ (.A1(_01582_),
    .A2(_01583_),
    .B1(_01584_),
    .B2(_01367_),
    .C(_01585_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06383_ (.I(_01564_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06384_ (.A1(net133),
    .A2(_01587_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06385_ (.I(net11),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06386_ (.I(_01589_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06387_ (.A1(_01586_),
    .A2(_01588_),
    .B(_01590_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06388_ (.I(_01324_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06389_ (.I(_01591_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06390_ (.A1(_01582_),
    .A2(\wb_counter[5] ),
    .B1(_01584_),
    .B2(_01592_),
    .C(_01585_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06391_ (.A1(net134),
    .A2(_01587_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06392_ (.A1(_01593_),
    .A2(_01594_),
    .B(_01590_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06393_ (.A1(_01582_),
    .A2(\wb_counter[6] ),
    .B1(_01584_),
    .B2(_01320_),
    .C(_01585_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06394_ (.A1(net135),
    .A2(_01587_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06395_ (.A1(_01595_),
    .A2(_01596_),
    .B(_01590_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06396_ (.A1(_01582_),
    .A2(\wb_counter[7] ),
    .B1(_01584_),
    .B2(_01327_),
    .C(_01585_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06397_ (.A1(net136),
    .A2(_01587_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06398_ (.A1(_01597_),
    .A2(_01598_),
    .B(_01590_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06399_ (.I(_01548_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06400_ (.I(\as2650.debug_psu[0] ),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06401_ (.I(_01600_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06402_ (.I(_01559_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06403_ (.A1(_01599_),
    .A2(\wb_counter[8] ),
    .B1(_01601_),
    .B2(_01570_),
    .C(_01602_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06404_ (.I(_01564_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06405_ (.A1(net137),
    .A2(_01604_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06406_ (.I(_01589_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06407_ (.A1(_01603_),
    .A2(_01605_),
    .B(_01606_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06408_ (.I(\as2650.debug_psu[1] ),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06409_ (.I(_01607_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06410_ (.I(_01608_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06411_ (.I(_01552_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06412_ (.A1(_01599_),
    .A2(\wb_counter[9] ),
    .B1(_01609_),
    .B2(_01610_),
    .C(_01602_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06413_ (.A1(net138),
    .A2(_01604_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06414_ (.A1(_01611_),
    .A2(_01612_),
    .B(_01606_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06415_ (.I(\as2650.debug_psu[2] ),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06416_ (.I(_01613_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06417_ (.I(_01614_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06418_ (.A1(_01599_),
    .A2(\wb_counter[10] ),
    .B1(_01615_),
    .B2(_01610_),
    .C(_01602_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06419_ (.A1(net108),
    .A2(_01604_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06420_ (.A1(_01616_),
    .A2(_01617_),
    .B(_01606_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06421_ (.I(\as2650.debug_psu[3] ),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06422_ (.I(_01618_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06423_ (.A1(_01599_),
    .A2(\wb_counter[11] ),
    .B1(_01619_),
    .B2(_01610_),
    .C(_01602_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06424_ (.A1(net109),
    .A2(_01604_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06425_ (.A1(_01620_),
    .A2(_01621_),
    .B(_01606_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06426_ (.I(_01548_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06427_ (.I(\as2650.debug_psu[4] ),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06428_ (.I(_01559_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06429_ (.A1(_01622_),
    .A2(\wb_counter[12] ),
    .B1(_01623_),
    .B2(_01610_),
    .C(_01624_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06430_ (.I(_01564_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06431_ (.A1(net110),
    .A2(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06432_ (.I(_01589_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06433_ (.A1(_01625_),
    .A2(_01627_),
    .B(_01628_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06434_ (.I(\as2650.debug_psu[5] ),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06435_ (.I(_01629_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06436_ (.A1(_01622_),
    .A2(\wb_counter[13] ),
    .B1(_01630_),
    .B2(_01553_),
    .C(_01624_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06437_ (.A1(net111),
    .A2(_01626_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06438_ (.A1(_01631_),
    .A2(_01632_),
    .B(_01628_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06439_ (.I(net144),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06440_ (.A1(_01622_),
    .A2(\wb_counter[14] ),
    .B1(_01633_),
    .B2(_01553_),
    .C(_01624_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06441_ (.A1(net112),
    .A2(_01626_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06442_ (.A1(_01634_),
    .A2(_01635_),
    .B(_01628_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06443_ (.I(\as2650.debug_psu[7] ),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06444_ (.A1(_01622_),
    .A2(\wb_counter[15] ),
    .B1(_01636_),
    .B2(_01553_),
    .C(_01624_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06445_ (.A1(net113),
    .A2(_01626_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06446_ (.A1(_01637_),
    .A2(_01638_),
    .B(_01628_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06447_ (.I(_01547_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06448_ (.I(_01639_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06449_ (.I(_01551_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06450_ (.I(_01641_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06451_ (.I(_01559_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06452_ (.I(_01643_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06453_ (.A1(_01640_),
    .A2(\wb_counter[16] ),
    .B(_01642_),
    .C(_01644_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06454_ (.I(_01563_),
    .Z(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06455_ (.I(_01646_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06456_ (.A1(net114),
    .A2(_01647_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06457_ (.I(_01589_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06458_ (.A1(_01645_),
    .A2(_01648_),
    .B(_01649_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06459_ (.A1(_01640_),
    .A2(\wb_counter[17] ),
    .B(_01642_),
    .C(_01644_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06460_ (.A1(net115),
    .A2(_01647_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06461_ (.A1(_01650_),
    .A2(_01651_),
    .B(_01649_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06462_ (.A1(_01640_),
    .A2(\wb_counter[18] ),
    .B(_01642_),
    .C(_01644_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06463_ (.A1(net116),
    .A2(_01647_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06464_ (.A1(_01652_),
    .A2(_01653_),
    .B(_01649_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06465_ (.A1(_01640_),
    .A2(\wb_counter[19] ),
    .B(_01642_),
    .C(_01644_),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06466_ (.A1(net117),
    .A2(_01647_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06467_ (.A1(_01654_),
    .A2(_01655_),
    .B(_01649_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06468_ (.I(_01639_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06469_ (.I(_01641_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06470_ (.I(_01643_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06471_ (.A1(_01656_),
    .A2(\wb_counter[20] ),
    .B(_01657_),
    .C(_01658_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06472_ (.I(_01646_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06473_ (.A1(net119),
    .A2(_01660_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06474_ (.I(net11),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06475_ (.I(_01662_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06476_ (.A1(_01659_),
    .A2(_01661_),
    .B(_01663_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06477_ (.A1(_01656_),
    .A2(\wb_counter[21] ),
    .B(_01657_),
    .C(_01658_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06478_ (.A1(net120),
    .A2(_01660_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06479_ (.A1(_01664_),
    .A2(_01665_),
    .B(_01663_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06480_ (.A1(_01656_),
    .A2(\wb_counter[22] ),
    .B(_01657_),
    .C(_01658_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06481_ (.A1(net121),
    .A2(_01660_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06482_ (.A1(_01666_),
    .A2(_01667_),
    .B(_01663_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06483_ (.A1(_01656_),
    .A2(\wb_counter[23] ),
    .B(_01657_),
    .C(_01658_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06484_ (.A1(net122),
    .A2(_01660_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06485_ (.A1(_01668_),
    .A2(_01669_),
    .B(_01663_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06486_ (.I(_01639_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06487_ (.I(_01641_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06488_ (.I(_01560_),
    .Z(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06489_ (.A1(_01670_),
    .A2(\wb_counter[24] ),
    .B(_01671_),
    .C(_01672_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06490_ (.I(_01646_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06491_ (.A1(net123),
    .A2(_01674_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06492_ (.I(_01662_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06493_ (.A1(_01673_),
    .A2(_01675_),
    .B(_01676_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06494_ (.A1(_01670_),
    .A2(\wb_counter[25] ),
    .B(_01671_),
    .C(_01672_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06495_ (.A1(net124),
    .A2(_01674_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06496_ (.A1(_01677_),
    .A2(_01678_),
    .B(_01676_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06497_ (.A1(_01670_),
    .A2(\wb_counter[26] ),
    .B(_01671_),
    .C(_01672_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06498_ (.A1(net125),
    .A2(_01674_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06499_ (.A1(_01679_),
    .A2(_01680_),
    .B(_01676_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06500_ (.A1(_01670_),
    .A2(\wb_counter[27] ),
    .B(_01671_),
    .C(_01672_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06501_ (.A1(net126),
    .A2(_01674_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06502_ (.A1(_01681_),
    .A2(_01682_),
    .B(_01676_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06503_ (.I(_01639_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06504_ (.I(_01641_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06505_ (.I(_01560_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06506_ (.A1(_01683_),
    .A2(\wb_counter[28] ),
    .B(_01684_),
    .C(_01685_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06507_ (.I(_01646_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06508_ (.A1(net127),
    .A2(_01687_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06509_ (.I(_01662_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06510_ (.A1(_01686_),
    .A2(_01688_),
    .B(_01689_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06511_ (.A1(_01683_),
    .A2(\wb_counter[29] ),
    .B(_01684_),
    .C(_01685_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06512_ (.A1(net128),
    .A2(_01687_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06513_ (.A1(_01690_),
    .A2(_01691_),
    .B(_01689_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06514_ (.A1(_01683_),
    .A2(\wb_counter[30] ),
    .B(_01684_),
    .C(_01685_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06515_ (.A1(net130),
    .A2(_01687_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06516_ (.A1(_01692_),
    .A2(_01693_),
    .B(_01689_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06517_ (.A1(_01683_),
    .A2(\wb_counter[31] ),
    .B(_01684_),
    .C(_01685_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06518_ (.A1(net131),
    .A2(_01687_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06519_ (.A1(_01694_),
    .A2(_01695_),
    .B(_01689_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06520_ (.A1(_01545_),
    .A2(net380),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06521_ (.A1(net12),
    .A2(_01547_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06522_ (.A1(net48),
    .A2(_01696_),
    .A3(_01643_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06523_ (.A1(wb_debug_cc),
    .A2(_01697_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06524_ (.A1(net48),
    .A2(_01696_),
    .A3(_01643_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06525_ (.A1(net15),
    .A2(_01699_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06526_ (.I(_01662_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06527_ (.A1(_01698_),
    .A2(net342),
    .B(_01701_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06528_ (.A1(_01317_),
    .A2(net376),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06529_ (.A1(net26),
    .A2(_01699_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06530_ (.A1(_01702_),
    .A2(_01703_),
    .B(_01701_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06531_ (.A1(\web_behavior[0] ),
    .A2(_01697_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06532_ (.A1(net37),
    .A2(_01699_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06533_ (.A1(_01704_),
    .A2(net331),
    .B(_01701_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06534_ (.A1(\web_behavior[1] ),
    .A2(_01697_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06535_ (.A1(net40),
    .A2(_01699_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06536_ (.A1(_01706_),
    .A2(net308),
    .B(_01701_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06537_ (.A1(net48),
    .A2(net13),
    .A3(_01558_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06538_ (.I(_01708_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06539_ (.I(_01709_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06540_ (.I(_01708_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06541_ (.I(_01711_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06542_ (.I(_00502_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06543_ (.I(_01713_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06544_ (.A1(net15),
    .A2(_01712_),
    .B(_01714_),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06545_ (.A1(_01550_),
    .A2(_01710_),
    .B(_01715_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06546_ (.A1(_01550_),
    .A2(\wb_counter[1] ),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06547_ (.A1(net26),
    .A2(_01712_),
    .B(_01714_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06548_ (.A1(_01710_),
    .A2(_01716_),
    .B(net366),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06549_ (.A1(_01550_),
    .A2(\wb_counter[1] ),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06550_ (.A1(\wb_counter[2] ),
    .A2(_01718_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06551_ (.A1(net37),
    .A2(_01712_),
    .B(_01714_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06552_ (.A1(_01710_),
    .A2(_01719_),
    .B(_01720_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06553_ (.I(_01709_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06554_ (.A1(\wb_counter[0] ),
    .A2(\wb_counter[1] ),
    .A3(\wb_counter[2] ),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06555_ (.A1(\wb_counter[3] ),
    .A2(_01722_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06556_ (.A1(net40),
    .A2(_01709_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06557_ (.A1(_01721_),
    .A2(_01723_),
    .B(net391),
    .C(_01545_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06558_ (.I(\wb_counter[3] ),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06559_ (.A1(_01725_),
    .A2(_01722_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06560_ (.A1(_01583_),
    .A2(_01726_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06561_ (.A1(net304),
    .A2(_01712_),
    .B(_01714_),
    .ZN(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06562_ (.A1(_01710_),
    .A2(_01727_),
    .B(net305),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06563_ (.I(_01708_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06564_ (.I(_01729_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06565_ (.I(_01730_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06566_ (.A1(_01583_),
    .A2(_01726_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06567_ (.A1(\wb_counter[5] ),
    .A2(_01732_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06568_ (.I(_01711_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06569_ (.I(_01713_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06570_ (.A1(net272),
    .A2(_01734_),
    .B(_01735_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06571_ (.A1(_01731_),
    .A2(_01733_),
    .B(net273),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06572_ (.A1(_01583_),
    .A2(\wb_counter[5] ),
    .A3(_01726_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06573_ (.A1(\wb_counter[6] ),
    .A2(_01737_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06574_ (.A1(net268),
    .A2(_01734_),
    .B(_01735_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06575_ (.A1(_01731_),
    .A2(_01738_),
    .B(net269),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06576_ (.A1(\wb_counter[4] ),
    .A2(\wb_counter[5] ),
    .A3(\wb_counter[6] ),
    .A4(_01726_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06577_ (.A1(\wb_counter[7] ),
    .A2(_01740_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06578_ (.A1(net264),
    .A2(_01734_),
    .B(_01735_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06579_ (.A1(_01731_),
    .A2(_01741_),
    .B(net265),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06580_ (.I(\wb_counter[7] ),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06581_ (.A1(_01743_),
    .A2(_01740_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06582_ (.A1(\wb_counter[8] ),
    .A2(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06583_ (.A1(net284),
    .A2(_01734_),
    .B(_01735_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06584_ (.A1(_01731_),
    .A2(_01745_),
    .B(net285),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06585_ (.I(_01708_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06586_ (.I(_01747_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06587_ (.A1(\wb_counter[8] ),
    .A2(_01744_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06588_ (.A1(\wb_counter[9] ),
    .A2(_01749_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06589_ (.I(_01711_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06590_ (.I(_01713_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06591_ (.A1(net338),
    .A2(_01751_),
    .B(_01752_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06592_ (.A1(_01748_),
    .A2(_01750_),
    .B(net339),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06593_ (.A1(\wb_counter[9] ),
    .A2(_01749_),
    .B(\wb_counter[10] ),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06594_ (.A1(\wb_counter[9] ),
    .A2(\wb_counter[10] ),
    .A3(_01749_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06595_ (.A1(_01754_),
    .A2(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06596_ (.A1(net288),
    .A2(_01751_),
    .B(_01752_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06597_ (.A1(_01748_),
    .A2(_01756_),
    .B(net289),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06598_ (.A1(\wb_counter[11] ),
    .A2(_01755_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06599_ (.A1(net276),
    .A2(_01751_),
    .B(_01752_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06600_ (.A1(_01748_),
    .A2(_01758_),
    .B(net277),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06601_ (.A1(\wb_counter[11] ),
    .A2(_01755_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06602_ (.A1(\wb_counter[12] ),
    .A2(_01760_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06603_ (.A1(net280),
    .A2(_01751_),
    .B(_01752_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06604_ (.A1(_01748_),
    .A2(_01761_),
    .B(net281),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06605_ (.I(_01747_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06606_ (.A1(\wb_counter[11] ),
    .A2(\wb_counter[12] ),
    .A3(_01755_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06607_ (.A1(\wb_counter[13] ),
    .A2(_01764_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06608_ (.I(_01711_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06609_ (.I(_01713_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06610_ (.A1(net19),
    .A2(_01766_),
    .B(_01767_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06611_ (.A1(_01763_),
    .A2(_01765_),
    .B(net372),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06612_ (.I(\wb_counter[13] ),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06613_ (.A1(_01769_),
    .A2(_01764_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06614_ (.A1(\wb_counter[14] ),
    .A2(_01770_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06615_ (.A1(net20),
    .A2(_01766_),
    .B(_01767_),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06616_ (.A1(_01763_),
    .A2(_01771_),
    .B(net363),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06617_ (.A1(\wb_counter[14] ),
    .A2(_01770_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06618_ (.A1(\wb_counter[15] ),
    .A2(_01773_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06619_ (.A1(net21),
    .A2(_01766_),
    .B(_01767_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06620_ (.A1(_01763_),
    .A2(_01774_),
    .B(net348),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06621_ (.A1(\wb_counter[14] ),
    .A2(\wb_counter[15] ),
    .A3(_01770_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06622_ (.A1(\wb_counter[16] ),
    .A2(_01776_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06623_ (.A1(net22),
    .A2(_01766_),
    .B(_01767_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06624_ (.A1(_01763_),
    .A2(_01777_),
    .B(net357),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06625_ (.I(_01747_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06626_ (.I(\wb_counter[16] ),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06627_ (.A1(_01780_),
    .A2(_01776_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06628_ (.A1(\wb_counter[17] ),
    .A2(_01781_),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06629_ (.I(_01729_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06630_ (.I(_00502_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06631_ (.I(_01784_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06632_ (.A1(net23),
    .A2(_01783_),
    .B(_01785_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06633_ (.A1(_01779_),
    .A2(_01782_),
    .B(_01786_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06634_ (.A1(\wb_counter[17] ),
    .A2(_01781_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06635_ (.A1(\wb_counter[18] ),
    .A2(_01787_),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06636_ (.A1(net24),
    .A2(_01783_),
    .B(_01785_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06637_ (.A1(_01779_),
    .A2(_01788_),
    .B(net369),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06638_ (.A1(\wb_counter[17] ),
    .A2(\wb_counter[18] ),
    .A3(_01781_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06639_ (.A1(\wb_counter[19] ),
    .A2(_01790_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06640_ (.A1(net25),
    .A2(_01783_),
    .B(_01785_),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06641_ (.A1(_01779_),
    .A2(_01791_),
    .B(net345),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06642_ (.I(\wb_counter[19] ),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06643_ (.A1(_01793_),
    .A2(_01790_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06644_ (.A1(\wb_counter[20] ),
    .A2(_01794_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06645_ (.A1(net27),
    .A2(_01783_),
    .B(_01785_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06646_ (.A1(_01779_),
    .A2(_01795_),
    .B(net354),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06647_ (.I(_01747_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06648_ (.A1(\wb_counter[20] ),
    .A2(_01794_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06649_ (.A1(\wb_counter[21] ),
    .A2(_01798_),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06650_ (.I(_01729_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06651_ (.I(_01784_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06652_ (.A1(net28),
    .A2(_01800_),
    .B(_01801_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06653_ (.A1(_01797_),
    .A2(_01799_),
    .B(net360),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06654_ (.A1(\wb_counter[20] ),
    .A2(\wb_counter[21] ),
    .A3(_01794_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06655_ (.A1(\wb_counter[22] ),
    .A2(_01803_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06656_ (.A1(net29),
    .A2(_01800_),
    .B(_01801_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06657_ (.A1(_01797_),
    .A2(_01804_),
    .B(net351),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06658_ (.I(\wb_counter[22] ),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06659_ (.A1(_01806_),
    .A2(_01803_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06660_ (.A1(\wb_counter[23] ),
    .A2(_01807_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06661_ (.A1(net296),
    .A2(_01800_),
    .B(_01801_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06662_ (.A1(_01797_),
    .A2(_01808_),
    .B(net297),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06663_ (.A1(\wb_counter[23] ),
    .A2(_01807_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06664_ (.A1(\wb_counter[24] ),
    .A2(_01810_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06665_ (.A1(net323),
    .A2(_01800_),
    .B(_01801_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06666_ (.A1(_01797_),
    .A2(_01811_),
    .B(net324),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06667_ (.I(_01709_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06668_ (.A1(\wb_counter[23] ),
    .A2(\wb_counter[24] ),
    .A3(_01807_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06669_ (.A1(\wb_counter[25] ),
    .A2(_01814_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06670_ (.I(_01729_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06671_ (.I(_01784_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06672_ (.A1(net319),
    .A2(_01816_),
    .B(_01817_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06673_ (.A1(_01813_),
    .A2(_01815_),
    .B(net320),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06674_ (.I(\wb_counter[25] ),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06675_ (.A1(_01819_),
    .A2(_01814_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06676_ (.A1(\wb_counter[26] ),
    .A2(_01820_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06677_ (.A1(net311),
    .A2(_01816_),
    .B(_01817_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06678_ (.A1(_01813_),
    .A2(_01821_),
    .B(net312),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06679_ (.A1(\wb_counter[26] ),
    .A2(_01820_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06680_ (.A1(\wb_counter[27] ),
    .A2(_01823_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06681_ (.A1(net300),
    .A2(_01816_),
    .B(_01817_),
    .ZN(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06682_ (.A1(_01813_),
    .A2(_01824_),
    .B(net301),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06683_ (.A1(\wb_counter[26] ),
    .A2(\wb_counter[27] ),
    .A3(_01820_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06684_ (.A1(\wb_counter[28] ),
    .A2(_01826_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06685_ (.A1(net315),
    .A2(_01816_),
    .B(_01817_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06686_ (.A1(_01813_),
    .A2(_01827_),
    .B(net316),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06687_ (.I(\wb_counter[28] ),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06688_ (.A1(_01829_),
    .A2(_01826_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06689_ (.A1(\wb_counter[29] ),
    .A2(_01830_),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06690_ (.I(_01784_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06691_ (.A1(net327),
    .A2(_01730_),
    .B(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06692_ (.A1(_01721_),
    .A2(_01831_),
    .B(net328),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06693_ (.A1(\wb_counter[29] ),
    .A2(_01830_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06694_ (.A1(\wb_counter[30] ),
    .A2(_01834_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06695_ (.A1(net292),
    .A2(_01730_),
    .B(_01832_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06696_ (.A1(_01721_),
    .A2(_01835_),
    .B(net293),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06697_ (.A1(\wb_counter[29] ),
    .A2(\wb_counter[30] ),
    .A3(_01830_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06698_ (.A1(\wb_counter[31] ),
    .A2(_01837_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06699_ (.A1(net334),
    .A2(_01730_),
    .B(_01832_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06700_ (.A1(_01721_),
    .A2(_01838_),
    .B(net335),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06701_ (.I(_01029_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06702_ (.I(\as2650.PC[0] ),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06703_ (.I(_01841_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06704_ (.A1(_01840_),
    .A2(_01842_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06705_ (.A1(_01034_),
    .A2(_01535_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06706_ (.A1(_00511_),
    .A2(_01844_),
    .B(_01178_),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06707_ (.A1(_01110_),
    .A2(_01129_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06708_ (.A1(_01189_),
    .A2(_01846_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06709_ (.I(_01847_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06710_ (.A1(_01068_),
    .A2(_01283_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06711_ (.A1(_01848_),
    .A2(_01849_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06712_ (.A1(_01055_),
    .A2(_01845_),
    .A3(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06713_ (.I(_01851_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06714_ (.I(_01852_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06715_ (.I(_01222_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06716_ (.I(_01112_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06717_ (.I(_01855_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06718_ (.A1(_01202_),
    .A2(_01393_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06719_ (.I(_00504_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06720_ (.A1(_01057_),
    .A2(_00956_),
    .A3(net232),
    .A4(_01044_),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06721_ (.I(_01859_),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06722_ (.A1(_01858_),
    .A2(_01860_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06723_ (.I(_01861_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06724_ (.I(_01862_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06725_ (.A1(_01857_),
    .A2(_01863_),
    .Z(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06726_ (.A1(_01856_),
    .A2(_01864_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06727_ (.I(_01865_),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06728_ (.I(_01866_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06729_ (.I(_01865_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06730_ (.I(_01868_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06731_ (.A1(_01556_),
    .A2(_01869_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06732_ (.I(_01851_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06733_ (.I(_01871_),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06734_ (.A1(_01854_),
    .A2(_01867_),
    .B(_01870_),
    .C(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06735_ (.A1(_01843_),
    .A2(_01853_),
    .B(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06736_ (.I(_01874_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06737_ (.A1(\as2650.debug_psu[2] ),
    .A2(\as2650.debug_psu[3] ),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06738_ (.I(\as2650.debug_psu[0] ),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06739_ (.A1(_01877_),
    .A2(_01607_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06740_ (.I(_01878_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06741_ (.I(_01879_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06742_ (.I(_01880_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06743_ (.I(_01881_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _06744_ (.A1(_01851_),
    .A2(_01864_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06745_ (.A1(_01882_),
    .A2(_01883_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06746_ (.A1(_01876_),
    .A2(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06747_ (.I(_01885_),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06748_ (.I(_01886_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06749_ (.I(_01885_),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06750_ (.A1(\as2650.stack[1][0] ),
    .A2(_01888_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06751_ (.A1(_01875_),
    .A2(_01887_),
    .B(_01889_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06752_ (.I(_01852_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06753_ (.I(_01840_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06754_ (.I(\as2650.PC[1] ),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06755_ (.I(_01892_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06756_ (.A1(_01842_),
    .A2(_01893_),
    .Z(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06757_ (.I(_01894_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06758_ (.A1(_01891_),
    .A2(_01893_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06759_ (.A1(_01891_),
    .A2(_01895_),
    .B(_01896_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06760_ (.I(_01442_),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06761_ (.I(_01868_),
    .Z(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06762_ (.A1(_01569_),
    .A2(_01899_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06763_ (.A1(_01898_),
    .A2(_01867_),
    .B(_01872_),
    .C(_01900_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06764_ (.A1(_01890_),
    .A2(_01897_),
    .B(_01901_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06765_ (.I(_01902_),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06766_ (.A1(\as2650.stack[1][1] ),
    .A2(_01888_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06767_ (.A1(_01887_),
    .A2(_01903_),
    .B(_01904_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06768_ (.I(_01029_),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06769_ (.I(_01905_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06770_ (.I(_01029_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06771_ (.A1(_01841_),
    .A2(_01892_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06772_ (.A1(_00571_),
    .A2(_01908_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06773_ (.I(_01909_),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06774_ (.I(_01910_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06775_ (.A1(_01907_),
    .A2(_01911_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06776_ (.A1(_01906_),
    .A2(_00571_),
    .B(_01912_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06777_ (.I(net251),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06778_ (.A1(_01574_),
    .A2(_01899_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06779_ (.A1(_01914_),
    .A2(_01867_),
    .B(_01872_),
    .C(_01915_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06780_ (.A1(_01890_),
    .A2(_01913_),
    .B(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06781_ (.I(_01917_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06782_ (.A1(\as2650.stack[1][2] ),
    .A2(_01888_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06783_ (.A1(_01887_),
    .A2(_01918_),
    .B(_01919_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06784_ (.I(_00562_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06785_ (.I(\as2650.PC[2] ),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06786_ (.A1(\as2650.PC[0] ),
    .A2(_01892_),
    .A3(_01921_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06787_ (.A1(_01920_),
    .A2(_01922_),
    .Z(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06788_ (.I(_01923_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06789_ (.I(_01924_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06790_ (.A1(_01907_),
    .A2(_01925_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06791_ (.A1(_01906_),
    .A2(_01920_),
    .B(_01926_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06792_ (.I(net386),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06793_ (.A1(_01579_),
    .A2(_01899_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06794_ (.A1(_01928_),
    .A2(_01867_),
    .B(_01872_),
    .C(_01929_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06795_ (.A1(_01890_),
    .A2(_01927_),
    .B(_01930_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06796_ (.I(_01931_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06797_ (.I(_01886_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06798_ (.A1(\as2650.stack[1][3] ),
    .A2(_01933_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06799_ (.A1(_01887_),
    .A2(_01932_),
    .B(_01934_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06800_ (.I(_01886_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06801_ (.I(_01935_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06802_ (.I(_01840_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06803_ (.I(_00575_),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06804_ (.I(_01840_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06805_ (.A1(_00562_),
    .A2(_01922_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06806_ (.A1(\as2650.PC[4] ),
    .A2(_01940_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06807_ (.I(_01941_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06808_ (.A1(_01939_),
    .A2(_01942_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06809_ (.A1(_01937_),
    .A2(_01938_),
    .B(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06810_ (.I(_01866_),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06811_ (.I(_01871_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06812_ (.I(_01358_),
    .Z(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06813_ (.I(_01947_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06814_ (.A1(_01948_),
    .A2(_01899_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06815_ (.A1(_01482_),
    .A2(_01945_),
    .B(_01946_),
    .C(_01949_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06816_ (.A1(_01890_),
    .A2(_01944_),
    .B(_01950_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06817_ (.I(_01951_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06818_ (.A1(\as2650.stack[1][4] ),
    .A2(_01933_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06819_ (.A1(_01936_),
    .A2(_01952_),
    .B(_01953_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06820_ (.I(_01852_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06821_ (.I(\as2650.PC[5] ),
    .Z(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06822_ (.A1(_00562_),
    .A2(_00575_),
    .A3(_01922_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06823_ (.A1(_01955_),
    .A2(_01956_),
    .Z(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06824_ (.I(_01957_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06825_ (.A1(_01939_),
    .A2(_01958_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06826_ (.A1(_01937_),
    .A2(_00560_),
    .B(_01959_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06827_ (.I(_01261_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06828_ (.I(_01961_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06829_ (.I(_01868_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06830_ (.A1(_01592_),
    .A2(_01963_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06831_ (.A1(_01962_),
    .A2(_01945_),
    .B(_01946_),
    .C(_01964_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06832_ (.A1(_01954_),
    .A2(_01960_),
    .B(_01965_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06833_ (.I(_01966_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06834_ (.A1(\as2650.stack[1][5] ),
    .A2(_01933_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06835_ (.A1(_01936_),
    .A2(_01967_),
    .B(_01968_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06836_ (.I(\as2650.PC[6] ),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06837_ (.A1(_01955_),
    .A2(_01956_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06838_ (.A1(_01969_),
    .A2(_01970_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06839_ (.I(_01971_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06840_ (.A1(_01907_),
    .A2(_01969_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06841_ (.A1(_01891_),
    .A2(_01972_),
    .B(_01973_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06842_ (.I(_01268_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06843_ (.A1(_01320_),
    .A2(_01963_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06844_ (.A1(_01975_),
    .A2(_01945_),
    .B(_01946_),
    .C(_01976_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06845_ (.A1(_01954_),
    .A2(_01974_),
    .B(_01977_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06846_ (.I(_01978_),
    .Z(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06847_ (.A1(\as2650.stack[1][6] ),
    .A2(_01933_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06848_ (.A1(_01936_),
    .A2(_01979_),
    .B(_01980_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06849_ (.I(\as2650.PC[7] ),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06850_ (.A1(\as2650.PC[5] ),
    .A2(_01969_),
    .A3(_01956_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06851_ (.A1(_01981_),
    .A2(_01982_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06852_ (.I(_01983_),
    .Z(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06853_ (.A1(_01907_),
    .A2(_01981_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06854_ (.A1(_01891_),
    .A2(_01984_),
    .B(_01985_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06855_ (.I(_01276_),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06856_ (.A1(_01327_),
    .A2(_01963_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06857_ (.A1(_01987_),
    .A2(_01945_),
    .B(_01946_),
    .C(_01988_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06858_ (.A1(_01954_),
    .A2(_01986_),
    .B(_01989_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06859_ (.I(_01990_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06860_ (.I(_01886_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06861_ (.A1(\as2650.stack[1][7] ),
    .A2(_01992_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06862_ (.A1(_01936_),
    .A2(_01991_),
    .B(_01993_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06863_ (.I(_01935_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06864_ (.I(\as2650.PC[8] ),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06865_ (.I(\as2650.PC[7] ),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06866_ (.A1(_01996_),
    .A2(_01982_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06867_ (.A1(_01995_),
    .A2(_01997_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06868_ (.I(_01998_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06869_ (.I(_01995_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06870_ (.I0(_01999_),
    .I1(_02000_),
    .S(_01905_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06871_ (.I(net104),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06872_ (.I(_01866_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06873_ (.I(_01871_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06874_ (.A1(_01600_),
    .A2(_01963_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06875_ (.A1(_02002_),
    .A2(_02003_),
    .B(_02004_),
    .C(_02005_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06876_ (.A1(_01954_),
    .A2(_02001_),
    .B(_02006_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06877_ (.I(_02007_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06878_ (.A1(\as2650.stack[1][8] ),
    .A2(_01992_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06879_ (.A1(_01994_),
    .A2(_02008_),
    .B(_02009_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06880_ (.I(_01852_),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06881_ (.A1(_01995_),
    .A2(_01997_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06882_ (.A1(\as2650.PC[9] ),
    .A2(_02011_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06883_ (.I(_02012_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06884_ (.I(\as2650.PC[9] ),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06885_ (.I0(_02013_),
    .I1(_02014_),
    .S(_01905_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06886_ (.I(net105),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06887_ (.I(_01868_),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06888_ (.A1(_01609_),
    .A2(_02017_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06889_ (.A1(_02016_),
    .A2(_02003_),
    .B(_02004_),
    .C(_02018_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06890_ (.A1(_02010_),
    .A2(_02015_),
    .B(_02019_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06891_ (.I(_02020_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06892_ (.A1(\as2650.stack[1][9] ),
    .A2(_01992_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06893_ (.A1(_01994_),
    .A2(_02021_),
    .B(_02022_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06894_ (.I(\as2650.PC[10] ),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06895_ (.I(_02023_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06896_ (.A1(_01995_),
    .A2(\as2650.PC[9] ),
    .A3(_01997_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06897_ (.A1(_02023_),
    .A2(_02025_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06898_ (.I(_02026_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06899_ (.I(_02027_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06900_ (.A1(_01939_),
    .A2(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06901_ (.A1(_01937_),
    .A2(_02024_),
    .B(_02029_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06902_ (.I(net74),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06903_ (.A1(_01614_),
    .A2(_02017_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06904_ (.A1(_02031_),
    .A2(_02003_),
    .B(_02004_),
    .C(_02032_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06905_ (.A1(_02010_),
    .A2(_02030_),
    .B(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06906_ (.I(_02034_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06907_ (.A1(\as2650.stack[1][10] ),
    .A2(_01992_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06908_ (.A1(_01994_),
    .A2(_02035_),
    .B(_02036_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06909_ (.I(\as2650.PC[11] ),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06910_ (.I(_02037_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06911_ (.A1(_02024_),
    .A2(_02025_),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06912_ (.A1(_02037_),
    .A2(_02039_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06913_ (.I(_02040_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06914_ (.A1(_01939_),
    .A2(_02041_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06915_ (.A1(_01937_),
    .A2(_02038_),
    .B(_02042_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06916_ (.I(net75),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06917_ (.A1(_01619_),
    .A2(_02017_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06918_ (.A1(_02044_),
    .A2(_02003_),
    .B(_02004_),
    .C(_02045_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06919_ (.A1(_02010_),
    .A2(_02043_),
    .B(_02046_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06920_ (.I(_02047_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06921_ (.A1(\as2650.stack[1][11] ),
    .A2(_01935_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06922_ (.A1(_01994_),
    .A2(_02048_),
    .B(_02049_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06923_ (.A1(_02037_),
    .A2(_02039_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06924_ (.A1(\as2650.PC[12] ),
    .A2(_02050_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06925_ (.I(\as2650.PC[12] ),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06926_ (.I0(_02051_),
    .I1(_02052_),
    .S(_01905_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06927_ (.I(net76),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06928_ (.I(_01866_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06929_ (.I(_01871_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06930_ (.A1(\as2650.debug_psu[4] ),
    .A2(_02017_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06931_ (.A1(_02054_),
    .A2(_02055_),
    .B(_02056_),
    .C(_02057_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06932_ (.A1(_02010_),
    .A2(_02053_),
    .B(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06933_ (.I(_02059_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06934_ (.A1(\as2650.stack[1][12] ),
    .A2(_01935_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06935_ (.A1(_01888_),
    .A2(_02060_),
    .B(_02061_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06936_ (.I(_01876_),
    .Z(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06937_ (.I(_01884_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06938_ (.A1(_02062_),
    .A2(_02063_),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06939_ (.I(_02064_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06940_ (.I(\as2650.page_reg[0] ),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06941_ (.I(_01332_),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06942_ (.A1(_01629_),
    .A2(_01869_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06943_ (.A1(_02067_),
    .A2(_02055_),
    .B(_02056_),
    .C(_02068_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06944_ (.A1(_02066_),
    .A2(_01853_),
    .B(_02069_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06945_ (.I(_02070_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06946_ (.A1(\as2650.stack[1][13] ),
    .A2(_02065_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06947_ (.A1(_02065_),
    .A2(_02071_),
    .B(_02072_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06948_ (.I(\as2650.page_reg[1] ),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06949_ (.I(_01342_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06950_ (.A1(net144),
    .A2(_01869_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06951_ (.A1(_02074_),
    .A2(_02055_),
    .B(_02056_),
    .C(_02075_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06952_ (.A1(_02073_),
    .A2(_01853_),
    .B(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06953_ (.I(_02077_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06954_ (.A1(\as2650.stack[1][14] ),
    .A2(_02064_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06955_ (.A1(_02065_),
    .A2(_02078_),
    .B(_02079_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06956_ (.I(_01355_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06957_ (.I(_02080_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06958_ (.A1(_01636_),
    .A2(_01869_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06959_ (.A1(_02081_),
    .A2(_02055_),
    .B(_02056_),
    .C(_02082_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06960_ (.A1(_00949_),
    .A2(_01853_),
    .B(_02083_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06961_ (.I(_02084_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06962_ (.A1(\as2650.stack[1][15] ),
    .A2(_02064_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06963_ (.A1(_02065_),
    .A2(_02085_),
    .B(_02086_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06964_ (.I(net6),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06965_ (.I(_02087_),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06966_ (.I(_02088_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06967_ (.I(_02089_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06968_ (.A1(\as2650.cycle[4] ),
    .A2(_01298_),
    .A3(_01284_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06969_ (.A1(_01054_),
    .A2(_02091_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06970_ (.I(_02092_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06971_ (.I(_02092_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06972_ (.A1(_01180_),
    .A2(_01471_),
    .A3(_01040_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06973_ (.I(_02095_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06974_ (.I(_02096_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06975_ (.A1(_01386_),
    .A2(_01422_),
    .A3(_01423_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06976_ (.A1(net6),
    .A2(_01153_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06977_ (.I(_02099_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06978_ (.A1(_02098_),
    .A2(_02100_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06979_ (.A1(\as2650.debug_psl[0] ),
    .A2(\as2650.debug_psl[3] ),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06980_ (.A1(_01386_),
    .A2(_01228_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06981_ (.A1(_01424_),
    .A2(_02099_),
    .A3(_02103_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06982_ (.A1(_01153_),
    .A2(_01422_),
    .A3(_01423_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06983_ (.A1(_02098_),
    .A2(_02100_),
    .B1(_02105_),
    .B2(_02103_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06984_ (.I(_02106_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06985_ (.A1(_02104_),
    .A2(_02107_),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06986_ (.A1(_02102_),
    .A2(_02108_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06987_ (.A1(_01118_),
    .A2(_01108_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06988_ (.A1(_01071_),
    .A2(_02110_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06989_ (.A1(_02102_),
    .A2(_02108_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06990_ (.A1(_02111_),
    .A2(_02112_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06991_ (.A1(_01383_),
    .A2(_02110_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06992_ (.A1(_01318_),
    .A2(\as2650.debug_psl[3] ),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06993_ (.A1(_02104_),
    .A2(_02106_),
    .B(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06994_ (.A1(_02108_),
    .A2(_02115_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06995_ (.A1(_02114_),
    .A2(_02116_),
    .A3(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06996_ (.A1(_01197_),
    .A2(_02107_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06997_ (.A1(_01113_),
    .A2(_02104_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06998_ (.A1(_01138_),
    .A2(_02107_),
    .B(_02119_),
    .C(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06999_ (.A1(_02109_),
    .A2(_02113_),
    .B(_02118_),
    .C(_02121_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07000_ (.A1(_01082_),
    .A2(_01118_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07001_ (.A1(_00612_),
    .A2(_02123_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07002_ (.I0(_02101_),
    .I1(_02122_),
    .S(_02124_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07003_ (.I(_02125_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07004_ (.A1(_01018_),
    .A2(_01083_),
    .A3(_01149_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07005_ (.A1(_01146_),
    .A2(_02127_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07006_ (.A1(_01855_),
    .A2(_01026_),
    .B(_01135_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07007_ (.A1(_01205_),
    .A2(_01288_),
    .A3(_02128_),
    .A4(_02129_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07008_ (.A1(_01531_),
    .A2(_01175_),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07009_ (.A1(_01054_),
    .A2(_02130_),
    .A3(_02131_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07010_ (.I(_02132_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07011_ (.I(_02133_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07012_ (.A1(_01089_),
    .A2(_01203_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07013_ (.A1(_01862_),
    .A2(_02135_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07014_ (.I(_02136_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07015_ (.I(_02137_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07016_ (.I(_01577_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07017_ (.I(_02102_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07018_ (.A1(_02139_),
    .A2(_00795_),
    .B(_02140_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07019_ (.I(_01438_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07020_ (.I(_01861_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07021_ (.A1(_01017_),
    .A2(_01209_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07022_ (.A1(_01383_),
    .A2(_01198_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07023_ (.A1(_02144_),
    .A2(_02145_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07024_ (.A1(_02143_),
    .A2(_02146_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07025_ (.I(_02147_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07026_ (.I(_02148_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07027_ (.A1(_01210_),
    .A2(_01287_),
    .A3(_02143_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07028_ (.I(_02150_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07029_ (.I(_00847_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07030_ (.A1(_01112_),
    .A2(_01390_),
    .A3(_02127_),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _07031_ (.A1(_00504_),
    .A2(_01859_),
    .A3(_02153_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07032_ (.I(_02154_),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07033_ (.I0(_02152_),
    .I1(_01102_),
    .S(_02155_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07034_ (.A1(_01136_),
    .A2(_01150_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07035_ (.A1(_01210_),
    .A2(_01287_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07036_ (.A1(_02157_),
    .A2(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07037_ (.A1(_01862_),
    .A2(_02159_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07038_ (.I(_02147_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07039_ (.A1(_01854_),
    .A2(_02151_),
    .B1(_02156_),
    .B2(_02160_),
    .C(_02161_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07040_ (.A1(_02142_),
    .A2(_02149_),
    .B(_02137_),
    .C(_02162_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07041_ (.A1(_02138_),
    .A2(_02141_),
    .B(_02163_),
    .C(_02133_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07042_ (.A1(_02126_),
    .A2(_02134_),
    .B(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07043_ (.A1(_02097_),
    .A2(_02165_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07044_ (.A1(_00825_),
    .A2(_02097_),
    .B(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07045_ (.A1(_02094_),
    .A2(_02167_),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07046_ (.A1(_02090_),
    .A2(_02093_),
    .B(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07047_ (.I(_02169_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07048_ (.A1(\as2650.insin[1] ),
    .A2(_01213_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07049_ (.A1(_02171_),
    .A2(_00662_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07050_ (.A1(\as2650.insin[0] ),
    .A2(_01213_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07051_ (.A1(_02173_),
    .A2(_00656_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07052_ (.A1(_02172_),
    .A2(_02174_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07053_ (.I(_02175_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07054_ (.I(_02172_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07055_ (.I(_02177_),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07056_ (.I(_01507_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07057_ (.I(_02128_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07058_ (.A1(_01205_),
    .A2(_01288_),
    .A3(_02180_),
    .A4(_02129_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07059_ (.I(_02181_),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07060_ (.A1(_01217_),
    .A2(_02182_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07061_ (.A1(_01180_),
    .A2(_02179_),
    .A3(_02183_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07062_ (.I(_02184_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07063_ (.I(_01121_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07064_ (.I(_02186_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07065_ (.I(_02187_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07066_ (.A1(_01359_),
    .A2(_02188_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07067_ (.A1(_02178_),
    .A2(_02185_),
    .A3(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07068_ (.I(_02190_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07069_ (.A1(_01321_),
    .A2(_01022_),
    .A3(_01533_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07070_ (.I(net381),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07071_ (.A1(_02193_),
    .A2(_01189_),
    .A3(_01109_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07072_ (.A1(_02192_),
    .A2(_02194_),
    .B(_01180_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07073_ (.A1(_01214_),
    .A2(_01167_),
    .A3(_01168_),
    .A4(_01038_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07074_ (.A1(_01053_),
    .A2(_02196_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07075_ (.I(_02197_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07076_ (.A1(_01115_),
    .A2(_01130_),
    .A3(_02198_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07077_ (.I(_02154_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07078_ (.A1(_02143_),
    .A2(_02159_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07079_ (.A1(_01145_),
    .A2(_02143_),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07080_ (.I(_02202_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07081_ (.A1(_02200_),
    .A2(_02201_),
    .A3(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07082_ (.A1(_02199_),
    .A2(_02204_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07083_ (.A1(_02148_),
    .A2(_02132_),
    .A3(_02092_),
    .A4(_02095_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07084_ (.A1(_02195_),
    .A2(_02137_),
    .A3(_02205_),
    .A4(_02206_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07085_ (.A1(_01359_),
    .A2(_02207_),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07086_ (.A1(_02176_),
    .A2(_02191_),
    .A3(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07087_ (.I(_02209_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07088_ (.I(_02126_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07089_ (.I(_02190_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07090_ (.I(_00650_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07091_ (.A1(_02148_),
    .A2(_02132_),
    .A3(_02203_),
    .A4(_02136_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07092_ (.A1(_01054_),
    .A2(_02091_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07093_ (.A1(_01507_),
    .A2(_01055_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07094_ (.A1(_02200_),
    .A2(_02201_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07095_ (.A1(_02199_),
    .A2(_02215_),
    .A3(_02216_),
    .A4(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _07096_ (.A1(_02195_),
    .A2(_02214_),
    .A3(_02218_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07097_ (.A1(_02213_),
    .A2(_02219_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07098_ (.I(_02220_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07099_ (.I(_00506_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07100_ (.A1(_02176_),
    .A2(_02221_),
    .B(_02190_),
    .C(_02222_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07101_ (.I(_02223_),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07102_ (.A1(_02211_),
    .A2(_02212_),
    .B1(_02224_),
    .B2(\as2650.regs[7][0] ),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07103_ (.A1(_02170_),
    .A2(_02210_),
    .B(_02225_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07104_ (.I(net7),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07105_ (.I(_02226_),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07106_ (.I(_02227_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07107_ (.I(_02228_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07108_ (.I(_02094_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07109_ (.I(_02134_),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07110_ (.A1(_01425_),
    .A2(_02100_),
    .A3(_02103_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07111_ (.A1(_01445_),
    .A2(_01447_),
    .B(_01387_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07112_ (.A1(net7),
    .A2(_01153_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07113_ (.I(_02234_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07114_ (.A1(_01445_),
    .A2(_01447_),
    .B(_01154_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07115_ (.I(_01385_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07116_ (.A1(_02237_),
    .A2(_01236_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07117_ (.A1(_02233_),
    .A2(_02235_),
    .B1(_02236_),
    .B2(_02238_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07118_ (.A1(_01448_),
    .A2(_02235_),
    .A3(_02238_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07119_ (.A1(_02239_),
    .A2(_02240_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07120_ (.A1(_02140_),
    .A2(_02232_),
    .B(_02107_),
    .C(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07121_ (.A1(_02140_),
    .A2(_02232_),
    .B(_02106_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07122_ (.A1(_02239_),
    .A2(_02240_),
    .A3(_02243_),
    .B(_02111_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07123_ (.I(_02123_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07124_ (.A1(_00612_),
    .A2(_02245_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07125_ (.A1(_02233_),
    .A2(_02235_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07126_ (.A1(_02105_),
    .A2(_02103_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07127_ (.A1(_02098_),
    .A2(_02100_),
    .A3(_02248_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07128_ (.A1(_02116_),
    .A2(_02241_),
    .A3(_02249_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07129_ (.A1(_01200_),
    .A2(_00840_),
    .B(_01443_),
    .C(_01440_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07130_ (.A1(_01460_),
    .A2(_01438_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07131_ (.I(_01152_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07132_ (.A1(_02251_),
    .A2(_02252_),
    .B(_02253_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07133_ (.I(_02234_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07134_ (.A1(_02251_),
    .A2(_02252_),
    .B(_02237_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07135_ (.A1(_02253_),
    .A2(_01442_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _07136_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02256_),
    .B2(_02257_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07137_ (.A1(_01448_),
    .A2(_02235_),
    .A3(_02238_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07138_ (.A1(_02258_),
    .A2(_02259_),
    .B1(_02249_),
    .B2(_02116_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07139_ (.A1(_01140_),
    .A2(_02260_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07140_ (.A1(_01148_),
    .A2(_02258_),
    .B(_02259_),
    .C(_01063_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07141_ (.A1(_01383_),
    .A2(_02258_),
    .B(_02262_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07142_ (.A1(_02246_),
    .A2(_02247_),
    .B1(_02250_),
    .B2(_02261_),
    .C(_02263_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07143_ (.A1(_02242_),
    .A2(_02244_),
    .B(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07144_ (.I(_02265_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07145_ (.I(_02134_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07146_ (.I(_02136_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07147_ (.I(_02268_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07148_ (.I(_02161_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07149_ (.I(_02268_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07150_ (.I(_02202_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07151_ (.I(_02272_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07152_ (.A1(_01591_),
    .A2(_01434_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07153_ (.I(_02150_),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07154_ (.I(_02155_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07155_ (.I(_02201_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07156_ (.I(_02155_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07157_ (.A1(_01105_),
    .A2(_02278_),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07158_ (.A1(_01434_),
    .A2(_02276_),
    .B(_02277_),
    .C(_02279_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07159_ (.I(_02203_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07160_ (.A1(_01898_),
    .A2(_02275_),
    .B(_02280_),
    .C(_02281_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07161_ (.I(_02161_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07162_ (.A1(_02273_),
    .A2(_02274_),
    .B(_02282_),
    .C(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07163_ (.A1(_01457_),
    .A2(_02270_),
    .B(_02271_),
    .C(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07164_ (.A1(_02152_),
    .A2(_02269_),
    .B(_02285_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07165_ (.A1(_02267_),
    .A2(_02286_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07166_ (.I(_02096_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07167_ (.A1(_02231_),
    .A2(_02266_),
    .B(_02287_),
    .C(_02288_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07168_ (.I(_02216_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07169_ (.I(_02215_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07170_ (.A1(_00840_),
    .A2(_02290_),
    .B(_02291_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07171_ (.A1(_02289_),
    .A2(_02292_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07172_ (.A1(_02229_),
    .A2(_02230_),
    .B(_02293_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07173_ (.I(_02223_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07174_ (.I(_02266_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07175_ (.I(_02190_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07176_ (.A1(\as2650.regs[7][1] ),
    .A2(_02295_),
    .B1(_02296_),
    .B2(_02297_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07177_ (.A1(_02210_),
    .A2(_02294_),
    .B(_02298_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07178_ (.I(net8),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07179_ (.I(_02299_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07180_ (.I(_02300_),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07181_ (.I(_02301_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07182_ (.I(_02124_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07183_ (.A1(_02237_),
    .A2(_01462_),
    .A3(_01463_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07184_ (.A1(net8),
    .A2(_02253_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07185_ (.A1(_02304_),
    .A2(_02305_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07186_ (.A1(_01154_),
    .A2(_01462_),
    .A3(_01463_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07187_ (.A1(_02237_),
    .A2(_01243_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07188_ (.A1(_02304_),
    .A2(_02305_),
    .B1(_02307_),
    .B2(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07189_ (.I(_02309_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07190_ (.I(_01386_),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07191_ (.A1(_00518_),
    .A2(_02311_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07192_ (.I(_02308_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07193_ (.A1(_01462_),
    .A2(_01463_),
    .B(_02312_),
    .C(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07194_ (.A1(_02310_),
    .A2(_02314_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07195_ (.A1(_02240_),
    .A2(_02243_),
    .B(_02258_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07196_ (.A1(_02315_),
    .A2(_02316_),
    .B(_01143_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07197_ (.A1(_02315_),
    .A2(_02316_),
    .B(_02317_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07198_ (.A1(_02236_),
    .A2(_02238_),
    .B(_02247_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07199_ (.A1(_02260_),
    .A2(_02319_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07200_ (.A1(_02315_),
    .A2(_02320_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07201_ (.A1(_01138_),
    .A2(_02310_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07202_ (.A1(_01328_),
    .A2(_02310_),
    .B(_02314_),
    .C(_01113_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07203_ (.A1(_02114_),
    .A2(_02321_),
    .B1(_02322_),
    .B2(_02323_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07204_ (.A1(_02303_),
    .A2(_02306_),
    .B(_02318_),
    .C(_02324_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07205_ (.I(_02325_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07206_ (.I(_00846_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07207_ (.A1(_01591_),
    .A2(_01433_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07208_ (.A1(_02327_),
    .A2(_02328_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07209_ (.A1(_01100_),
    .A2(_02278_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07210_ (.A1(_01457_),
    .A2(_02276_),
    .B(_02277_),
    .C(_02330_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07211_ (.A1(net251),
    .A2(_02275_),
    .B(_02331_),
    .C(_02281_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07212_ (.A1(_02273_),
    .A2(_02329_),
    .B(_02332_),
    .C(_02283_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07213_ (.A1(_01470_),
    .A2(_02270_),
    .B(_02271_),
    .C(_02333_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07214_ (.A1(_02142_),
    .A2(_02269_),
    .B(_02334_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07215_ (.A1(_02267_),
    .A2(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07216_ (.A1(_02231_),
    .A2(_02326_),
    .B(_02336_),
    .C(_02288_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07217_ (.A1(_00987_),
    .A2(_02290_),
    .B(_02291_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07218_ (.A1(_02337_),
    .A2(_02338_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07219_ (.A1(_02302_),
    .A2(_02230_),
    .B(_02339_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07220_ (.I(_02326_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07221_ (.A1(\as2650.regs[7][2] ),
    .A2(_02295_),
    .B1(_02341_),
    .B2(_02297_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07222_ (.A1(_02210_),
    .A2(_02340_),
    .B(_02342_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07223_ (.I(_02246_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07224_ (.A1(_01493_),
    .A2(_01093_),
    .B1(_01473_),
    .B2(_01474_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07225_ (.A1(_01023_),
    .A2(_01387_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07226_ (.A1(_01387_),
    .A2(_02344_),
    .B(_02345_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07227_ (.I(_02111_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07228_ (.I0(_01251_),
    .I1(_02344_),
    .S(_02253_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07229_ (.A1(_02346_),
    .A2(_02348_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07230_ (.A1(_01464_),
    .A2(_02305_),
    .A3(_02308_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07231_ (.A1(_02350_),
    .A2(_02316_),
    .B(_02309_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07232_ (.A1(_02349_),
    .A2(_02351_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07233_ (.A1(_02347_),
    .A2(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07234_ (.I(_02114_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _07235_ (.A1(_02310_),
    .A2(_02314_),
    .B1(_02319_),
    .B2(_02260_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07236_ (.A1(_01388_),
    .A2(_01464_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07237_ (.A1(_02356_),
    .A2(_02313_),
    .B(_02306_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07238_ (.A1(_02355_),
    .A2(_02357_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07239_ (.A1(_02349_),
    .A2(_02358_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07240_ (.I(net9),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07241_ (.I0(_02360_),
    .I1(_02344_),
    .S(_02311_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07242_ (.I(_02348_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07243_ (.A1(_02361_),
    .A2(_02362_),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07244_ (.A1(_01197_),
    .A2(_02361_),
    .A3(_02362_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07245_ (.A1(_02361_),
    .A2(_02362_),
    .B(_02364_),
    .C(_01298_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07246_ (.A1(_01384_),
    .A2(_02363_),
    .B(_02365_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07247_ (.A1(_02354_),
    .A2(_02359_),
    .B(_02366_),
    .C(_02246_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07248_ (.A1(_02343_),
    .A2(_02346_),
    .B1(_02353_),
    .B2(_02367_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07249_ (.I(_02368_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07250_ (.I(_02133_),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07251_ (.A1(_02142_),
    .A2(_02327_),
    .B(_01324_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07252_ (.A1(_01472_),
    .A2(_02371_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07253_ (.A1(_01095_),
    .A2(_02200_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07254_ (.A1(_01470_),
    .A2(_02278_),
    .B(_02277_),
    .C(_02373_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07255_ (.A1(_01928_),
    .A2(_02275_),
    .B(_02374_),
    .C(_02272_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07256_ (.A1(_02273_),
    .A2(_02372_),
    .B(_02375_),
    .C(_02149_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07257_ (.A1(_00893_),
    .A2(_02270_),
    .B(_02138_),
    .C(_02376_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07258_ (.A1(_02327_),
    .A2(_02269_),
    .B(_02377_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07259_ (.A1(_02370_),
    .A2(_02378_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07260_ (.A1(_02231_),
    .A2(_02369_),
    .B(_02379_),
    .C(_02288_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07261_ (.A1(_00871_),
    .A2(_02290_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07262_ (.A1(_02093_),
    .A2(_02380_),
    .A3(_02381_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07263_ (.I(_01023_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07264_ (.I(_02215_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07265_ (.A1(_02383_),
    .A2(_02384_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07266_ (.A1(_02382_),
    .A2(_02385_),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07267_ (.I(_02369_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07268_ (.A1(\as2650.regs[7][3] ),
    .A2(_02295_),
    .B1(_02387_),
    .B2(_02297_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07269_ (.A1(_02210_),
    .A2(_02386_),
    .B(_02388_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07270_ (.I(_02209_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07271_ (.I(net10),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07272_ (.I(_02390_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07273_ (.I(_02391_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07274_ (.A1(_02390_),
    .A2(_01154_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07275_ (.A1(_01155_),
    .A2(_01484_),
    .B(_02393_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07276_ (.I(_02394_),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07277_ (.I(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07278_ (.A1(_02311_),
    .A2(_01259_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07279_ (.A1(_02311_),
    .A2(_01485_),
    .B(_02397_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07280_ (.A1(_02394_),
    .A2(_02398_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07281_ (.I(_02399_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07282_ (.A1(_02349_),
    .A2(_02351_),
    .B(_02363_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07283_ (.A1(_02400_),
    .A2(_02401_),
    .B(_01144_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07284_ (.A1(_02400_),
    .A2(_02401_),
    .B(_02402_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07285_ (.I(_02398_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07286_ (.A1(_02395_),
    .A2(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07287_ (.A1(_02394_),
    .A2(_02398_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07288_ (.A1(_02346_),
    .A2(_02362_),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07289_ (.A1(_02361_),
    .A2(_02348_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07290_ (.A1(_02363_),
    .A2(_02408_),
    .B1(_02357_),
    .B2(_02355_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _07291_ (.A1(_02405_),
    .A2(_02406_),
    .B1(_02407_),
    .B2(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07292_ (.A1(_02409_),
    .A2(_02407_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07293_ (.A1(_02400_),
    .A2(_02411_),
    .B(_01140_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07294_ (.A1(_02395_),
    .A2(_02404_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07295_ (.A1(_01328_),
    .A2(_02406_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07296_ (.A1(_02395_),
    .A2(_02404_),
    .B(_02414_),
    .C(_01298_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07297_ (.A1(_01384_),
    .A2(_02413_),
    .B(_02415_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07298_ (.A1(_02410_),
    .A2(_02412_),
    .B(_02416_),
    .C(_02343_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07299_ (.A1(_02343_),
    .A2(_02396_),
    .B1(_02403_),
    .B2(_02417_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07300_ (.I(_02418_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07301_ (.I(_01096_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07302_ (.I0(_02420_),
    .I1(_01097_),
    .S(_02155_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07303_ (.A1(_01482_),
    .A2(_02151_),
    .B1(_02421_),
    .B2(_02160_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07304_ (.A1(_02161_),
    .A2(_02422_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07305_ (.A1(_01492_),
    .A2(_02149_),
    .B(_02268_),
    .C(_02423_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07306_ (.A1(_01472_),
    .A2(_02138_),
    .B(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07307_ (.A1(_02370_),
    .A2(_02425_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07308_ (.A1(_02370_),
    .A2(_02419_),
    .B(_02426_),
    .C(_02097_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07309_ (.A1(_00900_),
    .A2(_00901_),
    .A3(_02096_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07310_ (.A1(_02094_),
    .A2(_02427_),
    .A3(_02428_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07311_ (.A1(_02392_),
    .A2(_02093_),
    .B(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07312_ (.I(_02430_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07313_ (.I(_02419_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07314_ (.A1(\as2650.regs[7][4] ),
    .A2(_02295_),
    .B1(_02432_),
    .B2(_02297_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07315_ (.A1(_02389_),
    .A2(_02431_),
    .B(_02433_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07316_ (.I(net2),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07317_ (.I(_02434_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07318_ (.I(_02435_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07319_ (.I(_02436_),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07320_ (.I(_02343_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07321_ (.A1(_01080_),
    .A2(_01389_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07322_ (.A1(_01390_),
    .A2(_01496_),
    .B(_02439_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07323_ (.I0(_02434_),
    .I1(_01496_),
    .S(_01388_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07324_ (.I0(net101),
    .I1(_01496_),
    .S(_01155_),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07325_ (.A1(_02441_),
    .A2(_02442_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07326_ (.A1(_02441_),
    .A2(_02442_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07327_ (.A1(_02443_),
    .A2(_02444_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07328_ (.A1(_02396_),
    .A2(_02404_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07329_ (.A1(_02410_),
    .A2(_02445_),
    .A3(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07330_ (.A1(_02410_),
    .A2(_02446_),
    .B(_02445_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07331_ (.A1(_01141_),
    .A2(_02448_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07332_ (.A1(_02399_),
    .A2(_02401_),
    .B(_02406_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07333_ (.A1(_02445_),
    .A2(_02450_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07334_ (.A1(_01148_),
    .A2(_02443_),
    .B(_02444_),
    .C(_02245_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07335_ (.A1(_02145_),
    .A2(_02443_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07336_ (.A1(_02246_),
    .A2(_02453_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07337_ (.A1(_01144_),
    .A2(_02451_),
    .B(_02452_),
    .C(_02454_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07338_ (.A1(_02447_),
    .A2(_02449_),
    .B(_02455_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07339_ (.A1(_02438_),
    .A2(_02440_),
    .B(_02456_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07340_ (.I(_02457_),
    .Z(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07341_ (.I(_01087_),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07342_ (.A1(_01318_),
    .A2(_02459_),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07343_ (.A1(_01091_),
    .A2(_02278_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07344_ (.A1(_01492_),
    .A2(_02276_),
    .B(_02461_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07345_ (.A1(_01962_),
    .A2(_02275_),
    .B1(_02462_),
    .B2(_02160_),
    .C(_02281_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07346_ (.A1(_02273_),
    .A2(_02460_),
    .B(_02463_),
    .C(_02283_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07347_ (.A1(_01505_),
    .A2(_02270_),
    .B(_02271_),
    .C(_02464_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07348_ (.A1(_02420_),
    .A2(_02269_),
    .B(_02465_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07349_ (.A1(_02267_),
    .A2(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07350_ (.A1(_02231_),
    .A2(_02458_),
    .B(_02467_),
    .C(_02288_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07351_ (.A1(_00877_),
    .A2(_00883_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07352_ (.A1(_02469_),
    .A2(_02290_),
    .B(_02291_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07353_ (.A1(_02468_),
    .A2(_02470_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07354_ (.A1(_02437_),
    .A2(_02230_),
    .B(_02471_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07355_ (.I(_02458_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07356_ (.A1(\as2650.regs[7][5] ),
    .A2(_02224_),
    .B1(_02473_),
    .B2(_02212_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07357_ (.A1(_02389_),
    .A2(_02472_),
    .B(_02474_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07358_ (.A1(_01065_),
    .A2(_01390_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07359_ (.A1(_01391_),
    .A2(_01512_),
    .B(_02475_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07360_ (.I0(_01064_),
    .I1(_01512_),
    .S(_01388_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07361_ (.I0(_01272_),
    .I1(_01512_),
    .S(_01155_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07362_ (.A1(_02477_),
    .A2(_02478_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07363_ (.A1(_02477_),
    .A2(_02478_),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07364_ (.A1(_02479_),
    .A2(_02480_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07365_ (.A1(_02440_),
    .A2(_02442_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07366_ (.A1(_02448_),
    .A2(_02481_),
    .A3(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07367_ (.A1(_02448_),
    .A2(_02482_),
    .B(_02481_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07368_ (.A1(_02354_),
    .A2(_02484_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07369_ (.A1(_02483_),
    .A2(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07370_ (.I(_02444_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07371_ (.A1(_02443_),
    .A2(_02450_),
    .B(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07372_ (.A1(_02481_),
    .A2(_02488_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07373_ (.A1(_01144_),
    .A2(_02489_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07374_ (.A1(_01321_),
    .A2(_02479_),
    .B(_02480_),
    .C(_02245_),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07375_ (.A1(_02145_),
    .A2(_02479_),
    .B(_02491_),
    .C(_02303_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07376_ (.A1(_02486_),
    .A2(_02490_),
    .A3(_02492_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07377_ (.A1(_02438_),
    .A2(_02476_),
    .B(_02493_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07378_ (.A1(_01318_),
    .A2(_02459_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07379_ (.A1(_01504_),
    .A2(_02495_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07380_ (.A1(_02198_),
    .A2(_02153_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07381_ (.A1(_01086_),
    .A2(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07382_ (.A1(_01504_),
    .A2(_02276_),
    .B(_02277_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07383_ (.A1(_01975_),
    .A2(_02151_),
    .B1(_02498_),
    .B2(_02499_),
    .C(_02272_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07384_ (.A1(_02281_),
    .A2(_02496_),
    .B(_02500_),
    .C(_02149_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07385_ (.A1(_01517_),
    .A2(_02283_),
    .B(_02138_),
    .C(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07386_ (.A1(_02459_),
    .A2(_02271_),
    .B(_02502_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07387_ (.A1(_02370_),
    .A2(_02503_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07388_ (.A1(_02267_),
    .A2(_02494_),
    .B(_02504_),
    .C(_02097_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07389_ (.A1(_01509_),
    .A2(_02216_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07390_ (.A1(_02093_),
    .A2(_02505_),
    .A3(_02506_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07391_ (.I(_01065_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07392_ (.A1(_02508_),
    .A2(_02291_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07393_ (.A1(_02507_),
    .A2(_02509_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07394_ (.I(_02494_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07395_ (.A1(\as2650.regs[7][6] ),
    .A2(_02224_),
    .B1(_02511_),
    .B2(_02212_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07396_ (.A1(_02389_),
    .A2(_02510_),
    .B(_02512_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07397_ (.I(_00529_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07398_ (.I(_02513_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07399_ (.A1(_01156_),
    .A2(_01520_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07400_ (.A1(_00529_),
    .A2(_01156_),
    .B(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07401_ (.A1(_01389_),
    .A2(_01520_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07402_ (.A1(_01389_),
    .A2(_01279_),
    .B(_02517_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07403_ (.A1(_02516_),
    .A2(_02518_),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07404_ (.A1(_02516_),
    .A2(_02518_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07405_ (.I(_02520_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07406_ (.A1(_02476_),
    .A2(_02478_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07407_ (.A1(_02484_),
    .A2(_02519_),
    .A3(_02521_),
    .A4(_02522_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07408_ (.I(_02519_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07409_ (.A1(_02524_),
    .A2(_02521_),
    .B1(_02522_),
    .B2(_02484_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07410_ (.A1(_01141_),
    .A2(_02523_),
    .A3(_02525_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07411_ (.A1(_02519_),
    .A2(_02520_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07412_ (.A1(_02477_),
    .A2(_02478_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07413_ (.A1(_02528_),
    .A2(_02488_),
    .B(_02480_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07414_ (.A1(_02527_),
    .A2(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07415_ (.A1(_01321_),
    .A2(_02519_),
    .B(_02521_),
    .C(_02245_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07416_ (.A1(_02145_),
    .A2(_02524_),
    .B(_02531_),
    .C(_02303_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07417_ (.A1(_02347_),
    .A2(_02530_),
    .B(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07418_ (.A1(_02438_),
    .A2(_02516_),
    .B1(_02526_),
    .B2(_02533_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07419_ (.I(_02534_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07420_ (.A1(_01078_),
    .A2(_02497_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07421_ (.A1(_01517_),
    .A2(_02200_),
    .B(_02201_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07422_ (.A1(_01987_),
    .A2(_02151_),
    .B1(_02536_),
    .B2(_02537_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07423_ (.A1(_02459_),
    .A2(_00779_),
    .B(_01554_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07424_ (.A1(_01517_),
    .A2(_02539_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07425_ (.A1(_02203_),
    .A2(_02540_),
    .B(_02148_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07426_ (.A1(_02272_),
    .A2(_02538_),
    .B(_02541_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07427_ (.I(_02146_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07428_ (.A1(_01863_),
    .A2(_02543_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07429_ (.A1(_01577_),
    .A2(_02152_),
    .B(_02115_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07430_ (.A1(_02544_),
    .A2(_02545_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07431_ (.A1(_02137_),
    .A2(_02546_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07432_ (.A1(_01505_),
    .A2(_02268_),
    .B1(_02542_),
    .B2(_02547_),
    .C(_02133_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07433_ (.A1(_02134_),
    .A2(_02535_),
    .B(_02548_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07434_ (.I0(_00906_),
    .I1(_02549_),
    .S(_02096_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07435_ (.A1(_02092_),
    .A2(_02550_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07436_ (.A1(_02514_),
    .A2(_02094_),
    .B(_02551_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07437_ (.I(_02552_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07438_ (.I(_02535_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07439_ (.A1(\as2650.regs[7][7] ),
    .A2(_02224_),
    .B1(_02554_),
    .B2(_02212_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07440_ (.A1(_02389_),
    .A2(_02553_),
    .B(_02555_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07441_ (.I(\as2650.debug_psu[2] ),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07442_ (.I(_02556_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07443_ (.I(_01618_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07444_ (.A1(_02557_),
    .A2(_02558_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07445_ (.A1(_01884_),
    .A2(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07446_ (.I(_02560_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07447_ (.I(_02561_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07448_ (.I(_02562_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07449_ (.I(_02560_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07450_ (.A1(\as2650.stack[5][0] ),
    .A2(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07451_ (.A1(_01875_),
    .A2(_02563_),
    .B(_02565_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07452_ (.A1(\as2650.stack[5][1] ),
    .A2(_02564_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07453_ (.A1(_01903_),
    .A2(_02563_),
    .B(_02566_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(\as2650.stack[5][2] ),
    .A2(_02564_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07455_ (.A1(_01918_),
    .A2(_02563_),
    .B(_02567_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07456_ (.I(_02561_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07457_ (.A1(\as2650.stack[5][3] ),
    .A2(_02568_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07458_ (.A1(_01932_),
    .A2(_02563_),
    .B(_02569_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07459_ (.I(_02562_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07460_ (.A1(\as2650.stack[5][4] ),
    .A2(_02568_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07461_ (.A1(_01952_),
    .A2(_02570_),
    .B(_02571_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07462_ (.A1(\as2650.stack[5][5] ),
    .A2(_02568_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07463_ (.A1(_01967_),
    .A2(_02570_),
    .B(_02572_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07464_ (.A1(\as2650.stack[5][6] ),
    .A2(_02568_),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07465_ (.A1(_01979_),
    .A2(_02570_),
    .B(_02573_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07466_ (.I(_02561_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07467_ (.A1(\as2650.stack[5][7] ),
    .A2(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07468_ (.A1(_01991_),
    .A2(_02570_),
    .B(_02575_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07469_ (.I(_02561_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07470_ (.A1(\as2650.stack[5][8] ),
    .A2(_02574_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07471_ (.A1(_02008_),
    .A2(_02576_),
    .B(_02577_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07472_ (.A1(\as2650.stack[5][9] ),
    .A2(_02574_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07473_ (.A1(_02021_),
    .A2(_02576_),
    .B(_02578_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07474_ (.A1(\as2650.stack[5][10] ),
    .A2(_02574_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07475_ (.A1(_02035_),
    .A2(_02576_),
    .B(_02579_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07476_ (.A1(\as2650.stack[5][11] ),
    .A2(_02562_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07477_ (.A1(_02048_),
    .A2(_02576_),
    .B(_02580_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07478_ (.A1(\as2650.stack[5][12] ),
    .A2(_02562_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07479_ (.A1(_02060_),
    .A2(_02564_),
    .B(_02581_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07480_ (.A1(_02063_),
    .A2(_02559_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07481_ (.I(_02582_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07482_ (.A1(\as2650.stack[5][13] ),
    .A2(_02583_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07483_ (.A1(_02071_),
    .A2(_02583_),
    .B(_02584_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07484_ (.A1(\as2650.stack[5][14] ),
    .A2(_02582_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07485_ (.A1(_02078_),
    .A2(_02583_),
    .B(_02585_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07486_ (.A1(\as2650.stack[5][15] ),
    .A2(_02582_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07487_ (.A1(_02085_),
    .A2(_02583_),
    .B(_02586_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07488_ (.A1(\as2650.debug_psu[0] ),
    .A2(\as2650.debug_psu[1] ),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07489_ (.I(_02587_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07490_ (.I(_02588_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07491_ (.I(_02589_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07492_ (.I(_02590_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07493_ (.I(_02591_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07494_ (.I(_02592_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07495_ (.I(_02593_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07496_ (.A1(_01864_),
    .A2(_01851_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07497_ (.I(_01613_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07498_ (.I(\as2650.debug_psu[3] ),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07499_ (.A1(_02596_),
    .A2(_02597_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07500_ (.A1(_02595_),
    .A2(_02598_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07501_ (.A1(_02594_),
    .A2(_02599_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07502_ (.I(_02600_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07503_ (.I(_02601_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07504_ (.I(_02602_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07505_ (.I(_02600_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07506_ (.A1(\as2650.stack[4][0] ),
    .A2(_02604_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07507_ (.A1(_01875_),
    .A2(_02603_),
    .B(_02605_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07508_ (.A1(\as2650.stack[4][1] ),
    .A2(_02604_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07509_ (.A1(_01903_),
    .A2(_02603_),
    .B(_02606_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07510_ (.A1(\as2650.stack[4][2] ),
    .A2(_02604_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07511_ (.A1(_01918_),
    .A2(_02603_),
    .B(_02607_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07512_ (.I(_02601_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07513_ (.A1(\as2650.stack[4][3] ),
    .A2(_02608_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07514_ (.A1(_01932_),
    .A2(_02603_),
    .B(_02609_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07515_ (.I(_02602_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07516_ (.A1(\as2650.stack[4][4] ),
    .A2(_02608_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07517_ (.A1(_01952_),
    .A2(_02610_),
    .B(_02611_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07518_ (.A1(\as2650.stack[4][5] ),
    .A2(_02608_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07519_ (.A1(_01967_),
    .A2(_02610_),
    .B(_02612_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07520_ (.A1(\as2650.stack[4][6] ),
    .A2(_02608_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07521_ (.A1(_01979_),
    .A2(_02610_),
    .B(_02613_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07522_ (.I(_02601_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07523_ (.A1(\as2650.stack[4][7] ),
    .A2(_02614_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07524_ (.A1(_01991_),
    .A2(_02610_),
    .B(_02615_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07525_ (.I(_02601_),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07526_ (.A1(\as2650.stack[4][8] ),
    .A2(_02614_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07527_ (.A1(_02008_),
    .A2(_02616_),
    .B(_02617_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07528_ (.A1(\as2650.stack[4][9] ),
    .A2(_02614_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07529_ (.A1(_02021_),
    .A2(_02616_),
    .B(_02618_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07530_ (.A1(\as2650.stack[4][10] ),
    .A2(_02614_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07531_ (.A1(_02035_),
    .A2(_02616_),
    .B(_02619_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07532_ (.A1(\as2650.stack[4][11] ),
    .A2(_02602_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07533_ (.A1(_02048_),
    .A2(_02616_),
    .B(_02620_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07534_ (.A1(\as2650.stack[4][12] ),
    .A2(_02602_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07535_ (.A1(_02060_),
    .A2(_02604_),
    .B(_02621_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07536_ (.I(_01877_),
    .Z(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07537_ (.I(_01607_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07538_ (.I(_02623_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07539_ (.A1(_02622_),
    .A2(_02624_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07540_ (.I(_01883_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07541_ (.A1(_02626_),
    .A2(_02559_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07542_ (.A1(_02625_),
    .A2(_02627_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07543_ (.I(_02628_),
    .Z(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07544_ (.A1(\as2650.stack[4][13] ),
    .A2(_02629_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07545_ (.A1(_02071_),
    .A2(_02629_),
    .B(_02630_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07546_ (.A1(\as2650.stack[4][14] ),
    .A2(_02628_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07547_ (.A1(_02078_),
    .A2(_02629_),
    .B(_02631_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07548_ (.A1(\as2650.stack[4][15] ),
    .A2(_02628_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07549_ (.A1(_02085_),
    .A2(_02629_),
    .B(_02632_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07550_ (.A1(\as2650.debug_psu[0] ),
    .A2(_02623_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07551_ (.I(_02633_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07552_ (.I(_02634_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07553_ (.I(_02635_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07554_ (.I(_02636_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07555_ (.I(_02637_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07556_ (.I(_02638_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07557_ (.A1(_02062_),
    .A2(_02626_),
    .A3(_02639_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07558_ (.I(_02640_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07559_ (.I(_02641_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07560_ (.I(_02642_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07561_ (.I(_02640_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07562_ (.A1(\as2650.stack[2][0] ),
    .A2(_02644_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07563_ (.A1(_01875_),
    .A2(_02643_),
    .B(_02645_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07564_ (.A1(\as2650.stack[2][1] ),
    .A2(_02644_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07565_ (.A1(_01903_),
    .A2(_02643_),
    .B(_02646_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07566_ (.A1(\as2650.stack[2][2] ),
    .A2(_02644_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07567_ (.A1(_01918_),
    .A2(_02643_),
    .B(_02647_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07568_ (.I(_02641_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07569_ (.A1(\as2650.stack[2][3] ),
    .A2(_02648_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07570_ (.A1(_01932_),
    .A2(_02643_),
    .B(_02649_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07571_ (.I(_02642_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07572_ (.A1(\as2650.stack[2][4] ),
    .A2(_02648_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07573_ (.A1(_01952_),
    .A2(_02650_),
    .B(_02651_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07574_ (.A1(\as2650.stack[2][5] ),
    .A2(_02648_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07575_ (.A1(_01967_),
    .A2(_02650_),
    .B(_02652_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07576_ (.A1(\as2650.stack[2][6] ),
    .A2(_02648_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07577_ (.A1(_01979_),
    .A2(_02650_),
    .B(_02653_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07578_ (.I(_02641_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07579_ (.A1(\as2650.stack[2][7] ),
    .A2(_02654_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07580_ (.A1(_01991_),
    .A2(_02650_),
    .B(_02655_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07581_ (.I(_02641_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07582_ (.A1(\as2650.stack[2][8] ),
    .A2(_02654_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07583_ (.A1(_02008_),
    .A2(_02656_),
    .B(_02657_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07584_ (.A1(\as2650.stack[2][9] ),
    .A2(_02654_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07585_ (.A1(_02021_),
    .A2(_02656_),
    .B(_02658_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07586_ (.A1(\as2650.stack[2][10] ),
    .A2(_02654_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07587_ (.A1(_02035_),
    .A2(_02656_),
    .B(_02659_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07588_ (.A1(\as2650.stack[2][11] ),
    .A2(_02642_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07589_ (.A1(_02048_),
    .A2(_02656_),
    .B(_02660_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07590_ (.A1(\as2650.stack[2][12] ),
    .A2(_02642_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07591_ (.A1(_02060_),
    .A2(_02644_),
    .B(_02661_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07592_ (.A1(_02622_),
    .A2(_01609_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07593_ (.A1(_02062_),
    .A2(_02626_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07594_ (.A1(_02662_),
    .A2(_02663_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07595_ (.I(_02664_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07596_ (.A1(\as2650.stack[2][13] ),
    .A2(_02665_),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07597_ (.A1(_02071_),
    .A2(_02665_),
    .B(_02666_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07598_ (.A1(\as2650.stack[2][14] ),
    .A2(_02664_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07599_ (.A1(_02078_),
    .A2(_02665_),
    .B(_02667_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07600_ (.A1(\as2650.stack[2][15] ),
    .A2(_02664_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07601_ (.A1(_02085_),
    .A2(_02665_),
    .B(_02668_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07602_ (.I(_01874_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07603_ (.A1(_01877_),
    .A2(_02624_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07604_ (.I(_02670_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07605_ (.I(_02671_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07606_ (.I(_02672_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07607_ (.I(_02673_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07608_ (.I(_02674_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07609_ (.I(_02675_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07610_ (.A1(_01613_),
    .A2(_01618_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07611_ (.A1(_02595_),
    .A2(_02677_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07612_ (.A1(_02676_),
    .A2(_02678_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07613_ (.I(_02679_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07614_ (.I(_02680_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07615_ (.I(_02681_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07616_ (.I(_02679_),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07617_ (.A1(\as2650.stack[15][0] ),
    .A2(_02683_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07618_ (.A1(_02669_),
    .A2(_02682_),
    .B(_02684_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07619_ (.I(_01902_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07620_ (.A1(\as2650.stack[15][1] ),
    .A2(_02683_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07621_ (.A1(_02685_),
    .A2(_02682_),
    .B(_02686_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07622_ (.I(_01917_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07623_ (.A1(\as2650.stack[15][2] ),
    .A2(_02683_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07624_ (.A1(_02687_),
    .A2(_02682_),
    .B(_02688_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07625_ (.I(_01931_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07626_ (.I(_02680_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07627_ (.A1(\as2650.stack[15][3] ),
    .A2(_02690_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07628_ (.A1(_02689_),
    .A2(_02682_),
    .B(_02691_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07629_ (.I(_01951_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07630_ (.I(_02681_),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07631_ (.A1(\as2650.stack[15][4] ),
    .A2(_02690_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07632_ (.A1(_02692_),
    .A2(_02693_),
    .B(_02694_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07633_ (.I(_01966_),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07634_ (.A1(\as2650.stack[15][5] ),
    .A2(_02690_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07635_ (.A1(_02695_),
    .A2(_02693_),
    .B(_02696_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07636_ (.I(_01978_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07637_ (.A1(\as2650.stack[15][6] ),
    .A2(_02690_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07638_ (.A1(_02697_),
    .A2(_02693_),
    .B(_02698_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07639_ (.I(_01990_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07640_ (.I(_02680_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07641_ (.A1(\as2650.stack[15][7] ),
    .A2(_02700_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07642_ (.A1(_02699_),
    .A2(_02693_),
    .B(_02701_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07643_ (.I(_02007_),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07644_ (.I(_02680_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07645_ (.A1(\as2650.stack[15][8] ),
    .A2(_02700_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07646_ (.A1(_02702_),
    .A2(_02703_),
    .B(_02704_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07647_ (.I(_02020_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07648_ (.A1(\as2650.stack[15][9] ),
    .A2(_02700_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07649_ (.A1(_02705_),
    .A2(_02703_),
    .B(_02706_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07650_ (.I(_02034_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07651_ (.A1(\as2650.stack[15][10] ),
    .A2(_02700_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07652_ (.A1(_02707_),
    .A2(_02703_),
    .B(_02708_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07653_ (.I(_02047_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07654_ (.A1(\as2650.stack[15][11] ),
    .A2(_02681_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07655_ (.A1(_02709_),
    .A2(_02703_),
    .B(_02710_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07656_ (.I(_02059_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07657_ (.A1(\as2650.stack[15][12] ),
    .A2(_02681_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07658_ (.A1(_02711_),
    .A2(_02683_),
    .B(_02712_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07659_ (.I(_02070_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07660_ (.A1(_01600_),
    .A2(_01607_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07661_ (.I(_02714_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07662_ (.A1(_01615_),
    .A2(_01619_),
    .A3(_02626_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07663_ (.A1(_02715_),
    .A2(_02716_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07664_ (.I(_02717_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07665_ (.A1(\as2650.stack[15][13] ),
    .A2(_02718_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07666_ (.A1(_02713_),
    .A2(_02718_),
    .B(_02719_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07667_ (.I(_02077_),
    .Z(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07668_ (.A1(\as2650.stack[15][14] ),
    .A2(_02717_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07669_ (.A1(_02720_),
    .A2(_02718_),
    .B(_02721_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07670_ (.I(_02084_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07671_ (.A1(\as2650.stack[15][15] ),
    .A2(_02717_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07672_ (.A1(_02722_),
    .A2(_02718_),
    .B(_02723_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07673_ (.I(_02674_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07674_ (.A1(_02062_),
    .A2(_01883_),
    .A3(_02724_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07675_ (.I(_02725_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07676_ (.I(_02726_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07677_ (.I(_02727_),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07678_ (.I(_02725_),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07679_ (.A1(\as2650.stack[3][0] ),
    .A2(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07680_ (.A1(_02669_),
    .A2(_02728_),
    .B(_02730_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07681_ (.A1(\as2650.stack[3][1] ),
    .A2(_02729_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07682_ (.A1(_02685_),
    .A2(_02728_),
    .B(_02731_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07683_ (.A1(\as2650.stack[3][2] ),
    .A2(_02729_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07684_ (.A1(_02687_),
    .A2(_02728_),
    .B(_02732_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07685_ (.I(_02726_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07686_ (.A1(\as2650.stack[3][3] ),
    .A2(_02733_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07687_ (.A1(_02689_),
    .A2(_02728_),
    .B(_02734_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07688_ (.I(_02727_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07689_ (.A1(\as2650.stack[3][4] ),
    .A2(_02733_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07690_ (.A1(_02692_),
    .A2(_02735_),
    .B(_02736_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07691_ (.A1(\as2650.stack[3][5] ),
    .A2(_02733_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07692_ (.A1(_02695_),
    .A2(_02735_),
    .B(_02737_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07693_ (.A1(\as2650.stack[3][6] ),
    .A2(_02733_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07694_ (.A1(_02697_),
    .A2(_02735_),
    .B(_02738_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07695_ (.I(_02726_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07696_ (.A1(\as2650.stack[3][7] ),
    .A2(_02739_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07697_ (.A1(_02699_),
    .A2(_02735_),
    .B(_02740_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07698_ (.I(_02726_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07699_ (.A1(\as2650.stack[3][8] ),
    .A2(_02739_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07700_ (.A1(_02702_),
    .A2(_02741_),
    .B(_02742_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07701_ (.A1(\as2650.stack[3][9] ),
    .A2(_02739_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07702_ (.A1(_02705_),
    .A2(_02741_),
    .B(_02743_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07703_ (.A1(\as2650.stack[3][10] ),
    .A2(_02739_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07704_ (.A1(_02707_),
    .A2(_02741_),
    .B(_02744_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07705_ (.A1(\as2650.stack[3][11] ),
    .A2(_02727_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07706_ (.A1(_02709_),
    .A2(_02741_),
    .B(_02745_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07707_ (.A1(\as2650.stack[3][12] ),
    .A2(_02727_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07708_ (.A1(_02711_),
    .A2(_02729_),
    .B(_02746_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07709_ (.A1(_02663_),
    .A2(_02715_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07710_ (.I(_02747_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07711_ (.A1(\as2650.stack[3][13] ),
    .A2(_02748_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07712_ (.A1(_02713_),
    .A2(_02748_),
    .B(_02749_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07713_ (.A1(\as2650.stack[3][14] ),
    .A2(_02747_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07714_ (.A1(_02720_),
    .A2(_02748_),
    .B(_02750_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07715_ (.A1(\as2650.stack[3][15] ),
    .A2(_02747_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07716_ (.A1(_02722_),
    .A2(_02748_),
    .B(_02751_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07717_ (.A1(_00991_),
    .A2(_01430_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07718_ (.I(_01294_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07719_ (.A1(\as2650.last_addr[0] ),
    .A2(_02753_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07720_ (.A1(_02752_),
    .A2(_02754_),
    .B(_01163_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07721_ (.A1(\as2650.last_addr[1] ),
    .A2(_01313_),
    .B(_01454_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07722_ (.A1(_01304_),
    .A2(_02755_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07723_ (.A1(\as2650.last_addr[2] ),
    .A2(_01295_),
    .B(_01468_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07724_ (.A1(_01529_),
    .A2(_02756_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07725_ (.A1(\as2650.last_addr[3] ),
    .A2(_01313_),
    .B(_01479_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07726_ (.A1(_01304_),
    .A2(_02757_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07727_ (.A1(\as2650.last_addr[4] ),
    .A2(_02753_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07728_ (.A1(_01489_),
    .A2(_02758_),
    .B(_01163_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07729_ (.A1(\as2650.last_addr[5] ),
    .A2(_02753_),
    .B(_01501_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07730_ (.A1(_01304_),
    .A2(_02759_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07731_ (.A1(_01003_),
    .A2(_01430_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07732_ (.A1(\as2650.last_addr[6] ),
    .A2(_02753_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07733_ (.A1(_02760_),
    .A2(_02761_),
    .B(_01163_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07734_ (.I(_01303_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07735_ (.A1(_01010_),
    .A2(_01430_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07736_ (.A1(\as2650.last_addr[7] ),
    .A2(_01313_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07737_ (.A1(_02762_),
    .A2(_02763_),
    .A3(_02764_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07738_ (.A1(_02599_),
    .A2(_02639_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07739_ (.I(_02765_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07740_ (.I(_02766_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07741_ (.I(_02767_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07742_ (.I(_02765_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07743_ (.A1(\as2650.stack[6][0] ),
    .A2(_02769_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07744_ (.A1(_02669_),
    .A2(_02768_),
    .B(_02770_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07745_ (.A1(\as2650.stack[6][1] ),
    .A2(_02769_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07746_ (.A1(_02685_),
    .A2(_02768_),
    .B(_02771_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07747_ (.A1(\as2650.stack[6][2] ),
    .A2(_02769_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07748_ (.A1(_02687_),
    .A2(_02768_),
    .B(_02772_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07749_ (.I(_02766_),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07750_ (.A1(\as2650.stack[6][3] ),
    .A2(_02773_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07751_ (.A1(_02689_),
    .A2(_02768_),
    .B(_02774_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07752_ (.I(_02767_),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07753_ (.A1(\as2650.stack[6][4] ),
    .A2(_02773_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07754_ (.A1(_02692_),
    .A2(_02775_),
    .B(_02776_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07755_ (.A1(\as2650.stack[6][5] ),
    .A2(_02773_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07756_ (.A1(_02695_),
    .A2(_02775_),
    .B(_02777_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07757_ (.A1(\as2650.stack[6][6] ),
    .A2(_02773_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07758_ (.A1(_02697_),
    .A2(_02775_),
    .B(_02778_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07759_ (.I(_02766_),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07760_ (.A1(\as2650.stack[6][7] ),
    .A2(_02779_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07761_ (.A1(_02699_),
    .A2(_02775_),
    .B(_02780_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07762_ (.I(_02766_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07763_ (.A1(\as2650.stack[6][8] ),
    .A2(_02779_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07764_ (.A1(_02702_),
    .A2(_02781_),
    .B(_02782_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07765_ (.A1(\as2650.stack[6][9] ),
    .A2(_02779_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07766_ (.A1(_02705_),
    .A2(_02781_),
    .B(_02783_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07767_ (.A1(\as2650.stack[6][10] ),
    .A2(_02779_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07768_ (.A1(_02707_),
    .A2(_02781_),
    .B(_02784_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07769_ (.A1(\as2650.stack[6][11] ),
    .A2(_02767_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07770_ (.A1(_02709_),
    .A2(_02781_),
    .B(_02785_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07771_ (.A1(\as2650.stack[6][12] ),
    .A2(_02767_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07772_ (.A1(_02711_),
    .A2(_02769_),
    .B(_02786_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07773_ (.A1(_02627_),
    .A2(_02662_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07774_ (.I(_02787_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07775_ (.A1(\as2650.stack[6][13] ),
    .A2(_02788_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07776_ (.A1(_02713_),
    .A2(_02788_),
    .B(_02789_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07777_ (.A1(\as2650.stack[6][14] ),
    .A2(_02787_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07778_ (.A1(_02720_),
    .A2(_02788_),
    .B(_02790_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07779_ (.A1(\as2650.stack[6][15] ),
    .A2(_02787_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07780_ (.A1(_02722_),
    .A2(_02788_),
    .B(_02791_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07781_ (.A1(_01043_),
    .A2(_01027_),
    .A3(_01047_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07782_ (.A1(_01537_),
    .A2(_02792_),
    .B(_01533_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07783_ (.I(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07784_ (.A1(_01049_),
    .A2(_02794_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07785_ (.I(_02795_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07786_ (.I(_01540_),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07787_ (.A1(_02797_),
    .A2(_01176_),
    .A3(_01033_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07788_ (.I(_01841_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07789_ (.I(_02799_),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07790_ (.I(\as2650.instruction_args_latch[8] ),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07791_ (.A1(_02087_),
    .A2(_01858_),
    .A3(_01530_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07792_ (.A1(_02801_),
    .A2(_01174_),
    .B(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07793_ (.A1(_02800_),
    .A2(_02803_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07794_ (.A1(_00606_),
    .A2(_01118_),
    .A3(_02175_),
    .A4(_01115_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07795_ (.A1(_02805_),
    .A2(_01535_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07796_ (.I(_02806_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07797_ (.I(_02806_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07798_ (.A1(_02808_),
    .A2(_02804_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07799_ (.A1(_02090_),
    .A2(_02807_),
    .B(_02809_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07800_ (.A1(_01538_),
    .A2(_02804_),
    .B1(_02810_),
    .B2(_02792_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07801_ (.A1(_00566_),
    .A2(_01043_),
    .A3(_01048_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07802_ (.I(_02812_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07803_ (.A1(_01858_),
    .A2(_01045_),
    .B(\as2650.instruction_args_latch[0] ),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07804_ (.A1(_02087_),
    .A2(_01052_),
    .A3(net381),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07805_ (.A1(_02814_),
    .A2(_02815_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07806_ (.A1(_02193_),
    .A2(_01166_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07807_ (.I(_02817_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07808_ (.A1(_02798_),
    .A2(_02811_),
    .A3(_02813_),
    .B1(_02816_),
    .B2(_02818_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07809_ (.I(_00508_),
    .Z(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07810_ (.I(_02820_),
    .Z(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07811_ (.A1(_00826_),
    .A2(_02796_),
    .B(_02819_),
    .C(_02821_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07812_ (.I(\as2650.indirect_target[1] ),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07813_ (.I(_01186_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07814_ (.I(_02812_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07815_ (.I(_02793_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07816_ (.A1(_01048_),
    .A2(_01536_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07817_ (.I(_02826_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07818_ (.A1(_02799_),
    .A2(_01893_),
    .Z(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07819_ (.A1(_02801_),
    .A2(_01174_),
    .B(_02802_),
    .C(_02799_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07820_ (.A1(_00505_),
    .A2(_01531_),
    .B(\as2650.instruction_args_latch[9] ),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07821_ (.A1(_02226_),
    .A2(_01052_),
    .A3(_01539_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07822_ (.A1(_02830_),
    .A2(_02831_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07823_ (.A1(_02828_),
    .A2(_02829_),
    .A3(_02832_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07824_ (.I(_02226_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07825_ (.I(_02834_),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07826_ (.I(_02806_),
    .Z(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07827_ (.A1(_02836_),
    .A2(_02833_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07828_ (.A1(_02835_),
    .A2(_02808_),
    .B(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07829_ (.A1(_00521_),
    .A2(_01165_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07830_ (.I(_02839_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07831_ (.A1(_02827_),
    .A2(_02833_),
    .B1(_02838_),
    .B2(_02840_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07832_ (.I(_01533_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07833_ (.A1(_02822_),
    .A2(_02825_),
    .B1(_02841_),
    .B2(_02842_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07834_ (.A1(_01858_),
    .A2(_01045_),
    .B(\as2650.instruction_args_latch[1] ),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07835_ (.A1(_02226_),
    .A2(_01052_),
    .A3(_02193_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07836_ (.A1(_02844_),
    .A2(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07837_ (.A1(_02824_),
    .A2(_02843_),
    .B1(_02846_),
    .B2(_02818_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07838_ (.A1(_02822_),
    .A2(_02823_),
    .B(_02847_),
    .C(_02821_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07839_ (.I0(_02299_),
    .I1(\as2650.instruction_args_latch[10] ),
    .S(_01015_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07840_ (.I(_02848_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07841_ (.I(_02849_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07842_ (.A1(_01894_),
    .A2(_02830_),
    .A3(_02831_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07843_ (.A1(_02830_),
    .A2(_02831_),
    .B(_01894_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07844_ (.A1(_02829_),
    .A2(_02851_),
    .B(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07845_ (.A1(_01910_),
    .A2(_02850_),
    .A3(_02853_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07846_ (.A1(_01111_),
    .A2(_00521_),
    .A3(_01117_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07847_ (.I(_02855_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07848_ (.A1(_02856_),
    .A2(_02854_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07849_ (.A1(_02302_),
    .A2(_02856_),
    .B(_02857_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07850_ (.A1(_01538_),
    .A2(_02854_),
    .B1(_02858_),
    .B2(_02792_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07851_ (.A1(_02798_),
    .A2(_02813_),
    .A3(_02859_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07852_ (.I(_02817_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07853_ (.I0(_02299_),
    .I1(\as2650.instruction_args_latch[2] ),
    .S(_01171_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07854_ (.A1(_02861_),
    .A2(_02862_),
    .B(_01303_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07855_ (.A1(_00572_),
    .A2(_02796_),
    .B(_02860_),
    .C(_02863_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07856_ (.I(_01015_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07857_ (.A1(\as2650.instruction_args_latch[11] ),
    .A2(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07858_ (.A1(_02383_),
    .A2(_01174_),
    .B(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07859_ (.I(_02866_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07860_ (.A1(_01910_),
    .A2(_02849_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07861_ (.A1(_01910_),
    .A2(_02849_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07862_ (.A1(_02868_),
    .A2(_02853_),
    .B(_02869_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07863_ (.A1(_01924_),
    .A2(_02867_),
    .A3(_02870_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07864_ (.A1(_02806_),
    .A2(_02871_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07865_ (.A1(_02383_),
    .A2(_02836_),
    .B(_02872_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07866_ (.A1(_02827_),
    .A2(_02871_),
    .B1(_02873_),
    .B2(_02839_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07867_ (.A1(_00563_),
    .A2(_02825_),
    .B1(_02874_),
    .B2(_02842_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07868_ (.I0(_02360_),
    .I1(\as2650.instruction_args_latch[3] ),
    .S(_01170_),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07869_ (.A1(_02824_),
    .A2(_02875_),
    .B1(_02876_),
    .B2(_02818_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07870_ (.A1(_00563_),
    .A2(_02823_),
    .B(_02877_),
    .C(_02821_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07871_ (.A1(_01178_),
    .A2(_01166_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07872_ (.I0(_02390_),
    .I1(\as2650.instruction_args_latch[12] ),
    .S(_02864_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07873_ (.A1(_01941_),
    .A2(_02879_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07874_ (.I(_02880_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07875_ (.A1(_01923_),
    .A2(_02866_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07876_ (.A1(_01923_),
    .A2(_02866_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07877_ (.A1(_02882_),
    .A2(_02870_),
    .B(_02883_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07878_ (.A1(_02881_),
    .A2(_02884_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07879_ (.A1(_02836_),
    .A2(_02885_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07880_ (.A1(_02392_),
    .A2(_02807_),
    .B(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07881_ (.A1(_01538_),
    .A2(_02885_),
    .B1(_02887_),
    .B2(_02792_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07882_ (.A1(\as2650.indirect_target[4] ),
    .A2(_02794_),
    .B1(_02888_),
    .B2(_02798_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _07883_ (.I(_02390_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07884_ (.A1(\as2650.instruction_args_latch[4] ),
    .A2(_01171_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07885_ (.A1(_02890_),
    .A2(_01172_),
    .B(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07886_ (.A1(\as2650.indirect_target[4] ),
    .A2(_01164_),
    .B1(_02861_),
    .B2(_02892_),
    .C(_01303_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07887_ (.A1(_02878_),
    .A2(_02889_),
    .B(_02893_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07888_ (.I0(_02434_),
    .I1(_00536_),
    .S(_02864_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07889_ (.A1(_01957_),
    .A2(_02894_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07890_ (.A1(_01957_),
    .A2(_02894_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07891_ (.A1(_02895_),
    .A2(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07892_ (.A1(_01923_),
    .A2(_02866_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07893_ (.A1(_01909_),
    .A2(_02849_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07894_ (.I(_02087_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07895_ (.I0(_02900_),
    .I1(_02801_),
    .S(_02864_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07896_ (.I(\as2650.instruction_args_latch[9] ),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07897_ (.A1(_01053_),
    .A2(_01539_),
    .B(_02902_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07898_ (.A1(_02834_),
    .A2(_00505_),
    .A3(_01531_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07899_ (.A1(_02828_),
    .A2(_02903_),
    .A3(_02904_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07900_ (.A1(_02903_),
    .A2(_02904_),
    .B(_02828_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07901_ (.A1(_02799_),
    .A2(_02901_),
    .A3(_02905_),
    .B(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07902_ (.A1(_01909_),
    .A2(_02848_),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07903_ (.A1(_02899_),
    .A2(_02907_),
    .B(_02908_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07904_ (.A1(_01924_),
    .A2(_02867_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07905_ (.A1(_02898_),
    .A2(_02909_),
    .B(_02910_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07906_ (.A1(_01941_),
    .A2(_02879_),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07907_ (.A1(_02881_),
    .A2(_02911_),
    .B(_02912_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07908_ (.A1(_02897_),
    .A2(_02913_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07909_ (.I(_01080_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07910_ (.A1(_02836_),
    .A2(_02914_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07911_ (.A1(_02915_),
    .A2(_02808_),
    .B(_02916_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07912_ (.A1(_02826_),
    .A2(_02914_),
    .B1(_02917_),
    .B2(_02839_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07913_ (.A1(_00559_),
    .A2(_02825_),
    .B1(_02918_),
    .B2(_02842_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07914_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_01171_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07915_ (.A1(_01080_),
    .A2(_01172_),
    .B(_02920_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07916_ (.A1(_02824_),
    .A2(_02919_),
    .B1(_02921_),
    .B2(_02818_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07917_ (.A1(_00559_),
    .A2(_02823_),
    .B(_02922_),
    .C(_02821_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07918_ (.I(_02855_),
    .Z(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07919_ (.I0(_01064_),
    .I1(_00629_),
    .S(_01014_),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07920_ (.A1(_01971_),
    .A2(_02924_),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07921_ (.A1(_02881_),
    .A2(_02911_),
    .B(_02895_),
    .C(_02912_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07922_ (.A1(_02896_),
    .A2(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07923_ (.A1(_02925_),
    .A2(_02927_),
    .Z(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07924_ (.I(_01064_),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07925_ (.I(_02929_),
    .Z(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07926_ (.A1(_02930_),
    .A2(_02856_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07927_ (.A1(_02923_),
    .A2(_02928_),
    .B(_02931_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07928_ (.A1(_01537_),
    .A2(_02928_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07929_ (.A1(_02840_),
    .A2(_02932_),
    .B(_02933_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07930_ (.A1(_00552_),
    .A2(_02825_),
    .B1(_02934_),
    .B2(_02842_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07931_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_01172_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07932_ (.A1(_01065_),
    .A2(_01173_),
    .B(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07933_ (.A1(_02824_),
    .A2(_02935_),
    .B1(_02937_),
    .B2(_02817_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07934_ (.I(_00508_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07935_ (.I(_02939_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07936_ (.A1(_00552_),
    .A2(_02823_),
    .B(_02938_),
    .C(_02940_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07937_ (.I(_02924_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07938_ (.A1(_01983_),
    .A2(_02941_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07939_ (.I(_02941_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07940_ (.A1(_01971_),
    .A2(_02943_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07941_ (.A1(_02896_),
    .A2(_02925_),
    .A3(_02926_),
    .B(_02944_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07942_ (.A1(_02942_),
    .A2(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07943_ (.I(_02930_),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07944_ (.I0(_02947_),
    .I1(_02946_),
    .S(_02856_),
    .Z(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07945_ (.A1(_02827_),
    .A2(_02946_),
    .B1(_02948_),
    .B2(_02840_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07946_ (.A1(_01534_),
    .A2(_02949_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07947_ (.A1(\as2650.indirect_target[7] ),
    .A2(_02794_),
    .B(_02950_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07948_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_01173_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07949_ (.A1(_01061_),
    .A2(_01173_),
    .B(_02952_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07950_ (.I(_02953_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07951_ (.I(_01050_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07952_ (.A1(\as2650.indirect_target[7] ),
    .A2(_01041_),
    .B(_01183_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07953_ (.A1(_02878_),
    .A2(_02951_),
    .B1(_02954_),
    .B2(_02955_),
    .C(_02956_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07954_ (.A1(_01998_),
    .A2(_02941_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07955_ (.I(_02941_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07956_ (.A1(_01998_),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07957_ (.A1(_02957_),
    .A2(_02959_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07958_ (.A1(_02942_),
    .A2(_02925_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07959_ (.A1(_02897_),
    .A2(_02961_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07960_ (.I(_02894_),
    .Z(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07961_ (.A1(_01941_),
    .A2(_02879_),
    .B1(_02963_),
    .B2(_01957_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07962_ (.A1(_02964_),
    .A2(_02896_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07963_ (.A1(_01971_),
    .A2(_01983_),
    .B(_02943_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07964_ (.A1(_02961_),
    .A2(_02965_),
    .B(_02966_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _07965_ (.A1(_02880_),
    .A2(_02884_),
    .A3(_02962_),
    .B(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07966_ (.A1(_02960_),
    .A2(_02968_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07967_ (.A1(_02808_),
    .A2(_02969_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07968_ (.A1(_02931_),
    .A2(_02970_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07969_ (.A1(_02827_),
    .A2(_02969_),
    .B1(_02971_),
    .B2(_02840_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07970_ (.A1(_01534_),
    .A2(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07971_ (.A1(\as2650.indirect_target[8] ),
    .A2(_02794_),
    .B(_02973_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07972_ (.A1(\as2650.indirect_target[8] ),
    .A2(_01041_),
    .B(_01183_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07973_ (.A1(_02955_),
    .A2(_02901_),
    .B1(_02878_),
    .B2(_02974_),
    .C(_02975_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07974_ (.I(_01049_),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07975_ (.I(_02832_),
    .Z(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07976_ (.I(_02793_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07977_ (.A1(_02012_),
    .A2(_02943_),
    .Z(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07978_ (.A1(_01998_),
    .A2(_02958_),
    .Z(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07979_ (.A1(_02957_),
    .A2(net252),
    .B(_02980_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07980_ (.A1(_02979_),
    .A2(_02981_),
    .Z(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07981_ (.A1(_01117_),
    .A2(_02793_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07982_ (.A1(\as2650.indirect_target[9] ),
    .A2(_02978_),
    .B1(_02982_),
    .B2(_02983_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07983_ (.A1(_02813_),
    .A2(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07984_ (.A1(\as2650.indirect_target[9] ),
    .A2(_01305_),
    .B1(_02976_),
    .B2(_02977_),
    .C(_02985_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07985_ (.A1(_01529_),
    .A2(_02986_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07986_ (.I(_00507_),
    .Z(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07987_ (.I(_02987_),
    .Z(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07988_ (.I(_02983_),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07989_ (.A1(_02878_),
    .A2(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07990_ (.I(_02943_),
    .Z(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07991_ (.A1(_02026_),
    .A2(_02991_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07992_ (.I(_02958_),
    .Z(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07993_ (.A1(_02960_),
    .A2(_02979_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07994_ (.A1(_02012_),
    .A2(_02993_),
    .B1(_02968_),
    .B2(_02994_),
    .C(_02980_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07995_ (.A1(_02992_),
    .A2(_02995_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07996_ (.A1(_02990_),
    .A2(_02996_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07997_ (.A1(\as2650.indirect_target[10] ),
    .A2(_02796_),
    .B1(_02850_),
    .B2(_02976_),
    .C(_02997_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07998_ (.A1(_02988_),
    .A2(_02998_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07999_ (.I(_02867_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08000_ (.A1(_02027_),
    .A2(_02993_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08001_ (.A1(_02027_),
    .A2(_02993_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08002_ (.A1(_03000_),
    .A2(_02995_),
    .B(_03001_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _08003_ (.A1(_02040_),
    .A2(_02993_),
    .A3(_03002_),
    .Z(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08004_ (.A1(\as2650.indirect_target[11] ),
    .A2(_02978_),
    .B1(_02983_),
    .B2(_03003_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08005_ (.A1(_02813_),
    .A2(_03004_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08006_ (.A1(\as2650.indirect_target[11] ),
    .A2(_01305_),
    .B1(_02976_),
    .B2(_02999_),
    .C(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08007_ (.A1(_02988_),
    .A2(_03006_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08008_ (.I(_02879_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08009_ (.I(_02958_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08010_ (.A1(_02041_),
    .A2(_03008_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08011_ (.A1(_02028_),
    .A2(_02041_),
    .B(_03008_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08012_ (.A1(_02992_),
    .A2(_02995_),
    .A3(_03009_),
    .B(_03010_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08013_ (.A1(_02051_),
    .A2(_02991_),
    .A3(_03011_),
    .Z(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08014_ (.A1(_02990_),
    .A2(_03012_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08015_ (.A1(\as2650.indirect_target[12] ),
    .A2(_02795_),
    .B1(_03007_),
    .B2(_02976_),
    .C(_03013_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08016_ (.A1(_02988_),
    .A2(_03014_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08017_ (.I0(_02066_),
    .I1(_02963_),
    .S(_00614_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08018_ (.A1(\as2650.indirect_target[13] ),
    .A2(_02978_),
    .B1(_02989_),
    .B2(_02066_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08019_ (.A1(_01050_),
    .A2(_03016_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08020_ (.A1(_02955_),
    .A2(_03015_),
    .B(_03017_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08021_ (.A1(_02988_),
    .A2(_03018_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08022_ (.I(_02987_),
    .Z(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08023_ (.A1(\as2650.indirect_target[14] ),
    .A2(_02978_),
    .B1(_02989_),
    .B2(_02073_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08024_ (.A1(_01050_),
    .A2(_03020_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08025_ (.I(_02073_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08026_ (.A1(_01020_),
    .A2(_03008_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08027_ (.A1(_03022_),
    .A2(_01020_),
    .B(_02817_),
    .C(_03023_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08028_ (.A1(_03021_),
    .A2(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08029_ (.A1(_03019_),
    .A2(_03025_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08030_ (.A1(_02955_),
    .A2(_02989_),
    .B(_00949_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08031_ (.A1(\as2650.indirect_target[15] ),
    .A2(_02796_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08032_ (.I(_02820_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08033_ (.A1(_03026_),
    .A2(_03027_),
    .B(_03028_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08034_ (.A1(_00942_),
    .A2(_01185_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08035_ (.A1(_00509_),
    .A2(_03029_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08036_ (.A1(_01059_),
    .A2(_00628_),
    .B1(_00627_),
    .B2(_02861_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08037_ (.A1(_03030_),
    .A2(_03031_),
    .Z(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08038_ (.I(_03032_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08039_ (.A1(_01059_),
    .A2(_00626_),
    .B1(_00634_),
    .B2(_02861_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08040_ (.A1(_03030_),
    .A2(_03033_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08041_ (.I(_03034_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08042_ (.I(_01218_),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08043_ (.A1(_01906_),
    .A2(_01186_),
    .A3(_01845_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08044_ (.A1(_01214_),
    .A2(_01906_),
    .B1(_01166_),
    .B2(_03036_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08045_ (.A1(_03035_),
    .A2(_03037_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08046_ (.A1(_00942_),
    .A2(_01192_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08047_ (.I(_01860_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08048_ (.I(_03039_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08049_ (.A1(_01161_),
    .A2(_03040_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08050_ (.A1(_01147_),
    .A2(_03041_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08051_ (.A1(_01142_),
    .A2(_03041_),
    .B(_03042_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08052_ (.A1(_01164_),
    .A2(_03038_),
    .B(_03043_),
    .C(_02940_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08053_ (.A1(_01527_),
    .A2(_03041_),
    .B(net98),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08054_ (.A1(_03019_),
    .A2(_03044_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08055_ (.I(\as2650.warmup[1] ),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08056_ (.A1(_01832_),
    .A2(net1),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08057_ (.A1(\as2650.warmup[0] ),
    .A2(_03045_),
    .B(_03046_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08058_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08059_ (.A1(_03046_),
    .A2(_03047_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08060_ (.I(_02193_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08061_ (.I(_03048_),
    .Z(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08062_ (.I(_03049_),
    .Z(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08063_ (.A1(_01058_),
    .A2(_03048_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08064_ (.I(_03051_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08065_ (.A1(_02090_),
    .A2(_03050_),
    .B1(_03052_),
    .B2(\as2650.instruction_args_latch[0] ),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08066_ (.A1(_03035_),
    .A2(_03053_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08067_ (.A1(\as2650.instruction_args_latch[1] ),
    .A2(_03052_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08068_ (.I(_03049_),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08069_ (.A1(_02229_),
    .A2(_03055_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08070_ (.I(_01218_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08071_ (.A1(_03054_),
    .A2(_03056_),
    .B(_03057_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08072_ (.A1(_02302_),
    .A2(_03050_),
    .B1(_03052_),
    .B2(\as2650.instruction_args_latch[2] ),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08073_ (.A1(_03035_),
    .A2(_03058_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08074_ (.I(_01219_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08075_ (.I(_02360_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08076_ (.I(_03060_),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08077_ (.I(_03061_),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08078_ (.A1(_03062_),
    .A2(_03050_),
    .B1(_03052_),
    .B2(\as2650.instruction_args_latch[3] ),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08079_ (.A1(_03059_),
    .A2(_03063_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08080_ (.I(_02391_),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08081_ (.I(_03051_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08082_ (.A1(_03064_),
    .A2(_03050_),
    .B1(_03065_),
    .B2(\as2650.instruction_args_latch[4] ),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08083_ (.A1(_03059_),
    .A2(_03066_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08084_ (.I(_03048_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08085_ (.A1(_02437_),
    .A2(_03067_),
    .B1(_03065_),
    .B2(\as2650.instruction_args_latch[5] ),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08086_ (.A1(_03059_),
    .A2(_03068_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08087_ (.A1(_02947_),
    .A2(_03067_),
    .B1(_03065_),
    .B2(\as2650.instruction_args_latch[6] ),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08088_ (.A1(_03059_),
    .A2(_03069_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08089_ (.I(_01219_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08090_ (.I(_02514_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08091_ (.A1(_03071_),
    .A2(_03067_),
    .B1(_03065_),
    .B2(\as2650.instruction_args_latch[7] ),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08092_ (.A1(_03070_),
    .A2(_03072_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08093_ (.I(_01540_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08094_ (.I(_03073_),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08095_ (.A1(_02090_),
    .A2(_03074_),
    .B1(_01543_),
    .B2(\as2650.instruction_args_latch[8] ),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08096_ (.A1(_03070_),
    .A2(_03075_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08097_ (.I(_03073_),
    .Z(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08098_ (.A1(_02229_),
    .A2(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08099_ (.I(_01542_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(\as2650.instruction_args_latch[9] ),
    .A2(_03078_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08101_ (.A1(_03077_),
    .A2(_03079_),
    .B(_03057_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08102_ (.A1(_02302_),
    .A2(_03074_),
    .B1(_01543_),
    .B2(\as2650.instruction_args_latch[10] ),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08103_ (.A1(_03070_),
    .A2(_03080_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08104_ (.A1(_03062_),
    .A2(_03074_),
    .B1(_01543_),
    .B2(\as2650.instruction_args_latch[11] ),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08105_ (.A1(_03070_),
    .A2(_03081_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08106_ (.A1(_03064_),
    .A2(_03074_),
    .B1(_01542_),
    .B2(\as2650.instruction_args_latch[12] ),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08107_ (.A1(_01219_),
    .A2(_03082_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08108_ (.A1(_02437_),
    .A2(_03076_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08109_ (.A1(_00536_),
    .A2(_03078_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08110_ (.A1(_03083_),
    .A2(_03084_),
    .B(_03057_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08111_ (.A1(_00629_),
    .A2(_03078_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08112_ (.A1(_02947_),
    .A2(_03076_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08113_ (.A1(_03085_),
    .A2(_03086_),
    .B(_03057_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08114_ (.A1(_03071_),
    .A2(_03076_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08115_ (.A1(\as2650.instruction_args_latch[15] ),
    .A2(_03078_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08116_ (.A1(_03087_),
    .A2(_03088_),
    .B(_03035_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08117_ (.I(_01847_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08118_ (.A1(_01046_),
    .A2(_03089_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08119_ (.I(_03090_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08120_ (.I(_02803_),
    .Z(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08121_ (.A1(_00604_),
    .A2(_02805_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08122_ (.I(_03093_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08123_ (.I(_03094_),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08124_ (.A1(_03095_),
    .A2(net96),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _08125_ (.A1(_02937_),
    .A2(_03096_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08126_ (.I(_03094_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08127_ (.A1(_03098_),
    .A2(net93),
    .B(_02892_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08128_ (.A1(_03094_),
    .A2(net91),
    .B(_02862_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08129_ (.A1(_03093_),
    .A2(net89),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08130_ (.A1(_02814_),
    .A2(_02815_),
    .B(_03101_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08131_ (.A1(_03093_),
    .A2(net90),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08132_ (.A1(_02844_),
    .A2(_02845_),
    .A3(_03103_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08133_ (.A1(_02844_),
    .A2(_02845_),
    .B(_03103_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08134_ (.A1(_03102_),
    .A2(_03104_),
    .B(_03105_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08135_ (.A1(_03095_),
    .A2(net91),
    .A3(_02862_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08136_ (.A1(_03100_),
    .A2(_03106_),
    .B(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08137_ (.I(_02876_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08138_ (.A1(_03094_),
    .A2(net92),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08139_ (.A1(_03109_),
    .A2(_03110_),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08140_ (.A1(_03109_),
    .A2(_03110_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08141_ (.A1(_03108_),
    .A2(_03111_),
    .B(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08142_ (.A1(_03095_),
    .A2(net93),
    .A3(_02892_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08143_ (.I(_03114_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08144_ (.A1(_03099_),
    .A2(_03113_),
    .B(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _08145_ (.A1(_03095_),
    .A2(net94),
    .A3(_02921_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08146_ (.A1(_03098_),
    .A2(net94),
    .B(_02921_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08147_ (.A1(_03117_),
    .A2(_03118_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _08148_ (.I(_03119_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08149_ (.A1(_03116_),
    .A2(_03120_),
    .B(_03117_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08150_ (.A1(_03098_),
    .A2(net97),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08151_ (.A1(_02953_),
    .A2(_03122_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08152_ (.A1(_02954_),
    .A2(_03122_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08153_ (.A1(_02937_),
    .A2(_03096_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08154_ (.A1(_02954_),
    .A2(_03122_),
    .B(_03125_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08155_ (.A1(_03126_),
    .A2(_03124_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _08156_ (.A1(_03097_),
    .A2(_03121_),
    .A3(_03123_),
    .B(_03127_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _08157_ (.A1(_03092_),
    .A2(_02977_),
    .A3(_02850_),
    .A4(_03128_),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08158_ (.A1(_02867_),
    .A2(_03007_),
    .A3(_03129_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08159_ (.A1(_02963_),
    .A2(_03130_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08160_ (.A1(_01876_),
    .A2(_02587_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08161_ (.A1(_01613_),
    .A2(_02625_),
    .B(\as2650.debug_psu[3] ),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08162_ (.A1(_03132_),
    .A2(_03133_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08163_ (.I(_03134_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08164_ (.I(_03135_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08165_ (.I(_03136_),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08166_ (.I(_03137_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08167_ (.I(_03138_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08168_ (.A1(\as2650.debug_psu[2] ),
    .A2(_02587_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08169_ (.I(_03140_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08170_ (.I(_03141_),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08171_ (.I(_03142_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08172_ (.I(_03143_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08173_ (.I(_03144_),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08174_ (.I(_01882_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08175_ (.I(_02637_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08176_ (.A1(\as2650.stack[4][13] ),
    .A2(_03146_),
    .B1(_03147_),
    .B2(\as2650.stack[5][13] ),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08177_ (.I(_02592_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08178_ (.A1(\as2650.stack[7][13] ),
    .A2(_03149_),
    .B1(_02724_),
    .B2(\as2650.stack[6][13] ),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08179_ (.A1(_03145_),
    .A2(_03148_),
    .A3(_03150_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08180_ (.A1(_02556_),
    .A2(_02588_),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08181_ (.I(_03152_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08182_ (.I(_03153_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08183_ (.I(_03154_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08184_ (.I(_03155_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08185_ (.A1(\as2650.stack[0][13] ),
    .A2(_03146_),
    .B1(_03147_),
    .B2(\as2650.stack[1][13] ),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08186_ (.A1(\as2650.stack[3][13] ),
    .A2(_03149_),
    .B1(_02724_),
    .B2(\as2650.stack[2][13] ),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08187_ (.A1(_03156_),
    .A2(_03157_),
    .A3(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08188_ (.A1(_03151_),
    .A2(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08189_ (.A1(\as2650.stack[11][13] ),
    .A2(_03149_),
    .B1(_02724_),
    .B2(\as2650.stack[10][13] ),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08190_ (.I(_01882_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08191_ (.A1(\as2650.stack[8][13] ),
    .A2(_03162_),
    .B1(_02638_),
    .B2(\as2650.stack[9][13] ),
    .C(_03145_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08192_ (.A1(\as2650.stack[15][13] ),
    .A2(_02593_),
    .B1(_02675_),
    .B2(\as2650.stack[14][13] ),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08193_ (.A1(\as2650.stack[12][13] ),
    .A2(_03162_),
    .B1(_02638_),
    .B2(\as2650.stack[13][13] ),
    .C(_03156_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08194_ (.A1(_03161_),
    .A2(_03163_),
    .B1(_03164_),
    .B2(_03165_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08195_ (.A1(_03139_),
    .A2(_03166_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08196_ (.A1(_03139_),
    .A2(_03160_),
    .B(_03167_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08197_ (.I(_02196_),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08198_ (.I(_03169_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08199_ (.I(_03170_),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08200_ (.I(_01136_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08201_ (.A1(_01120_),
    .A2(_03172_),
    .Z(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08202_ (.A1(_01127_),
    .A2(_03173_),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08203_ (.I(_03174_),
    .Z(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08204_ (.I(_03175_),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08205_ (.A1(_03171_),
    .A2(_03176_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08206_ (.I0(_03168_),
    .I1(_02066_),
    .S(_03177_),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08207_ (.I(_01846_),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08208_ (.A1(\as2650.page_reg[0] ),
    .A2(_02923_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08209_ (.A1(_01022_),
    .A2(_03179_),
    .A3(_01534_),
    .A4(_03180_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08210_ (.I(_03090_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08211_ (.A1(_03178_),
    .A2(_03181_),
    .B(_03182_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08212_ (.A1(_03091_),
    .A2(_03131_),
    .B(_03183_),
    .C(_02940_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08213_ (.A1(_02999_),
    .A2(_03007_),
    .A3(_02963_),
    .A4(_03129_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08214_ (.A1(_03008_),
    .A2(_03184_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08215_ (.I(_01539_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08216_ (.I(_03186_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08217_ (.A1(_01034_),
    .A2(_01535_),
    .A3(_03089_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08218_ (.I(_03188_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08219_ (.I(_03189_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08220_ (.A1(_02073_),
    .A2(_03187_),
    .A3(_02923_),
    .A4(_03190_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08221_ (.I(_03090_),
    .Z(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08222_ (.I(_03188_),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08223_ (.A1(\as2650.stack[4][14] ),
    .A2(_03146_),
    .B1(_03147_),
    .B2(\as2650.stack[5][14] ),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08224_ (.A1(\as2650.stack[7][14] ),
    .A2(_02593_),
    .B1(_02675_),
    .B2(\as2650.stack[6][14] ),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08225_ (.A1(_03145_),
    .A2(_03194_),
    .A3(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08226_ (.A1(\as2650.stack[0][14] ),
    .A2(_03146_),
    .B1(_03147_),
    .B2(\as2650.stack[1][14] ),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08227_ (.A1(\as2650.stack[3][14] ),
    .A2(_02593_),
    .B1(_02675_),
    .B2(\as2650.stack[2][14] ),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08228_ (.A1(_03156_),
    .A2(_03197_),
    .A3(_03198_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08229_ (.A1(_03196_),
    .A2(_03199_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08230_ (.A1(\as2650.stack[11][14] ),
    .A2(_02592_),
    .B1(_02674_),
    .B2(\as2650.stack[10][14] ),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08231_ (.A1(\as2650.stack[8][14] ),
    .A2(_03162_),
    .B1(_02637_),
    .B2(\as2650.stack[9][14] ),
    .C(_03145_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08232_ (.A1(\as2650.stack[15][14] ),
    .A2(_02592_),
    .B1(_02674_),
    .B2(\as2650.stack[14][14] ),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08233_ (.A1(\as2650.stack[12][14] ),
    .A2(_03162_),
    .B1(_02638_),
    .B2(\as2650.stack[13][14] ),
    .C(_03155_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08234_ (.A1(_03201_),
    .A2(_03202_),
    .B1(_03203_),
    .B2(_03204_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08235_ (.A1(_03138_),
    .A2(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08236_ (.A1(_03139_),
    .A2(_03200_),
    .B(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08237_ (.A1(_03177_),
    .A2(_03207_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08238_ (.A1(_03022_),
    .A2(_03177_),
    .B1(_03193_),
    .B2(_03073_),
    .C(_03208_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08239_ (.A1(_03192_),
    .A2(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08240_ (.I(_02939_),
    .Z(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08241_ (.A1(_03091_),
    .A2(_03185_),
    .B1(_03191_),
    .B2(_03210_),
    .C(_03211_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08242_ (.A1(_00537_),
    .A2(_01016_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08243_ (.A1(_00950_),
    .A2(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08244_ (.A1(_02991_),
    .A2(_03184_),
    .B(_03213_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08245_ (.A1(_02991_),
    .A2(_03184_),
    .A3(_03213_),
    .B(_03182_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08246_ (.I(_03215_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08247_ (.I(_03186_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08248_ (.A1(_03217_),
    .A2(_02807_),
    .A3(_03190_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08249_ (.A1(\as2650.stack[4][15] ),
    .A2(_01882_),
    .B1(_02637_),
    .B2(\as2650.stack[5][15] ),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08250_ (.I(_02588_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08251_ (.I(_03220_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08252_ (.I(_03221_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08253_ (.I(_02670_),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08254_ (.I(_03223_),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08255_ (.I(_03224_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08256_ (.A1(\as2650.stack[7][15] ),
    .A2(_03222_),
    .B1(_03225_),
    .B2(\as2650.stack[6][15] ),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08257_ (.A1(_03144_),
    .A2(_03219_),
    .A3(_03226_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08258_ (.I(_01878_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08259_ (.I(_03228_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08260_ (.I(_03229_),
    .Z(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08261_ (.I(_03230_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08262_ (.I(_02633_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08263_ (.I(_03232_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08264_ (.I(_03233_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08265_ (.I(_03234_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08266_ (.A1(\as2650.stack[0][15] ),
    .A2(_03231_),
    .B1(_03235_),
    .B2(\as2650.stack[1][15] ),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08267_ (.A1(\as2650.stack[3][15] ),
    .A2(_03222_),
    .B1(_03225_),
    .B2(\as2650.stack[2][15] ),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08268_ (.A1(_03155_),
    .A2(_03236_),
    .A3(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08269_ (.A1(_03227_),
    .A2(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08270_ (.A1(\as2650.stack[11][15] ),
    .A2(_03222_),
    .B1(_03225_),
    .B2(\as2650.stack[10][15] ),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08271_ (.I(_03140_),
    .Z(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08272_ (.I(_03241_),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08273_ (.I(_03242_),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08274_ (.A1(\as2650.stack[8][15] ),
    .A2(_03231_),
    .B1(_03235_),
    .B2(\as2650.stack[9][15] ),
    .C(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08275_ (.A1(\as2650.stack[15][15] ),
    .A2(_03222_),
    .B1(_03225_),
    .B2(\as2650.stack[14][15] ),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08276_ (.I(_03152_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08277_ (.I(_03246_),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08278_ (.I(_03247_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08279_ (.A1(\as2650.stack[12][15] ),
    .A2(_03231_),
    .B1(_03235_),
    .B2(\as2650.stack[13][15] ),
    .C(_03248_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08280_ (.A1(_03240_),
    .A2(_03244_),
    .B1(_03245_),
    .B2(_03249_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08281_ (.A1(_03138_),
    .A2(_03250_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08282_ (.A1(_03138_),
    .A2(_03239_),
    .B(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08283_ (.I0(_03252_),
    .I1(_00949_),
    .S(_03177_),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08284_ (.A1(_03218_),
    .A2(_03253_),
    .B(_03182_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08285_ (.A1(_03214_),
    .A2(_03216_),
    .B(_03254_),
    .C(_02940_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08286_ (.I(_02900_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08287_ (.I(_03169_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08288_ (.I(_03256_),
    .Z(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08289_ (.I(_03257_),
    .Z(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08290_ (.I(_03258_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08291_ (.I(_03171_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08292_ (.I(_03260_),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08293_ (.I(_01183_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08294_ (.A1(\as2650.insin[0] ),
    .A2(_03261_),
    .B(_03262_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08295_ (.A1(_03255_),
    .A2(_03259_),
    .B(_03263_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08296_ (.A1(\as2650.insin[1] ),
    .A2(_03261_),
    .B(_03262_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08297_ (.A1(_02835_),
    .A2(_03259_),
    .B(_03264_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08298_ (.I(_00518_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08299_ (.A1(\as2650.insin[2] ),
    .A2(_03261_),
    .B(_03262_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08300_ (.A1(_03265_),
    .A2(_03259_),
    .B(_03266_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08301_ (.A1(\as2650.insin[3] ),
    .A2(_03261_),
    .B(_03262_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08302_ (.A1(_02383_),
    .A2(_03259_),
    .B(_03267_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08303_ (.I(_03258_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08304_ (.I(_03260_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08305_ (.I(_01302_),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08306_ (.A1(\as2650.insin[4] ),
    .A2(_03269_),
    .B(_03270_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08307_ (.A1(_02890_),
    .A2(_03268_),
    .B(_03271_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08308_ (.A1(\as2650.insin[5] ),
    .A2(_03269_),
    .B(_03270_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08309_ (.A1(_02915_),
    .A2(_03268_),
    .B(_03272_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08310_ (.A1(\as2650.insin[6] ),
    .A2(_03269_),
    .B(_03270_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08311_ (.A1(_02508_),
    .A2(_03268_),
    .B(_03273_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08312_ (.I(_01061_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08313_ (.A1(\as2650.insin[7] ),
    .A2(_03269_),
    .B(_03270_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08314_ (.A1(_03274_),
    .A2(_03268_),
    .B(_03275_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08315_ (.I(_01309_),
    .Z(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08316_ (.A1(\as2650.last_addr[8] ),
    .A2(_03276_),
    .B(_01417_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08317_ (.A1(_03019_),
    .A2(_03277_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08318_ (.A1(\as2650.last_addr[9] ),
    .A2(_01310_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08319_ (.A1(_02762_),
    .A2(_01451_),
    .A3(_03278_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08320_ (.A1(\as2650.last_addr[10] ),
    .A2(_03276_),
    .B(_01459_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08321_ (.A1(_03019_),
    .A2(_03279_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08322_ (.A1(\as2650.last_addr[11] ),
    .A2(_01310_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08323_ (.A1(_02762_),
    .A2(_01477_),
    .A3(_03280_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08324_ (.A1(\as2650.last_addr[12] ),
    .A2(_03276_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08325_ (.A1(_01487_),
    .A2(_03281_),
    .B(_03028_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08326_ (.A1(\as2650.last_addr[13] ),
    .A2(_01310_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08327_ (.A1(_02762_),
    .A2(_01499_),
    .A3(_03282_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08328_ (.A1(\as2650.last_addr[14] ),
    .A2(_01297_),
    .B(_01506_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08329_ (.A1(_00510_),
    .A2(_03283_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08330_ (.A1(\as2650.last_addr[15] ),
    .A2(_03276_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08331_ (.A1(_01308_),
    .A2(_01522_),
    .A3(_03284_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08332_ (.I(_00594_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08333_ (.I(_03285_),
    .Z(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08334_ (.I(_01848_),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08335_ (.A1(_03286_),
    .A2(_03287_),
    .B(_03048_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08336_ (.I(_03288_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08337_ (.I(_02800_),
    .Z(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08338_ (.I(_03285_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08339_ (.A1(_03290_),
    .A2(_03291_),
    .B(_03190_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08340_ (.A1(_01848_),
    .A2(_01844_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08341_ (.I(_03293_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08342_ (.I(_03294_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08343_ (.I(_03186_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08344_ (.A1(_02810_),
    .A2(_03295_),
    .B(_03296_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08345_ (.I(_00556_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08346_ (.I(_03298_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08347_ (.I(_03293_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08348_ (.A1(_03299_),
    .A2(_03300_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08349_ (.A1(_01127_),
    .A2(_03173_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08350_ (.I(_03302_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08351_ (.I(_03303_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08352_ (.I(_03136_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08353_ (.I(_01879_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08354_ (.I(_02634_),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08355_ (.A1(\as2650.stack[4][0] ),
    .A2(_03306_),
    .B1(_03307_),
    .B2(\as2650.stack[5][0] ),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08356_ (.I(_02589_),
    .Z(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08357_ (.I(_02671_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08358_ (.A1(\as2650.stack[7][0] ),
    .A2(_03309_),
    .B1(_03310_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08359_ (.A1(_03242_),
    .A2(_03308_),
    .A3(_03311_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08360_ (.I(_03246_),
    .Z(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08361_ (.A1(\as2650.stack[0][0] ),
    .A2(_01880_),
    .B1(_03307_),
    .B2(\as2650.stack[1][0] ),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08362_ (.A1(\as2650.stack[3][0] ),
    .A2(_03309_),
    .B1(_03310_),
    .B2(\as2650.stack[2][0] ),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08363_ (.A1(_03313_),
    .A2(_03314_),
    .A3(_03315_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08364_ (.A1(_03312_),
    .A2(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08365_ (.I(_03135_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08366_ (.I(_02588_),
    .Z(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08367_ (.I(_03319_),
    .Z(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08368_ (.I(_02670_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08369_ (.I(_03321_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08370_ (.A1(\as2650.stack[11][0] ),
    .A2(_03320_),
    .B1(_03322_),
    .B2(\as2650.stack[10][0] ),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08371_ (.I(_03228_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08372_ (.I(_03232_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08373_ (.A1(\as2650.stack[8][0] ),
    .A2(_03324_),
    .B1(_03325_),
    .B2(\as2650.stack[9][0] ),
    .C(_03241_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08374_ (.A1(\as2650.stack[15][0] ),
    .A2(_03320_),
    .B1(_03322_),
    .B2(\as2650.stack[14][0] ),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08375_ (.A1(\as2650.stack[12][0] ),
    .A2(_03324_),
    .B1(_03325_),
    .B2(\as2650.stack[13][0] ),
    .C(_03153_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08376_ (.A1(_03323_),
    .A2(_03326_),
    .B1(_03327_),
    .B2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08377_ (.A1(_03318_),
    .A2(_03329_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08378_ (.A1(_03305_),
    .A2(_03317_),
    .B(_03330_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08379_ (.A1(_03290_),
    .A2(_03304_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08380_ (.A1(_03304_),
    .A2(_03331_),
    .B(_03332_),
    .C(_01196_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08381_ (.A1(_01020_),
    .A2(_03179_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08382_ (.I(_03334_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08383_ (.A1(_01030_),
    .A2(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08384_ (.I(_01194_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08385_ (.I(_03337_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08386_ (.A1(_02800_),
    .A2(_03336_),
    .B(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08387_ (.A1(_03290_),
    .A2(_03336_),
    .B(_03339_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08388_ (.I(_01860_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08389_ (.I(_03341_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08390_ (.A1(_03333_),
    .A2(_03340_),
    .B(_03342_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08391_ (.A1(_03290_),
    .A2(_03040_),
    .B1(_03301_),
    .B2(_01541_),
    .C(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08392_ (.I(_03344_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08393_ (.A1(_03292_),
    .A2(_03297_),
    .B(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08394_ (.I(_00556_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08395_ (.I(_03347_),
    .Z(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08396_ (.A1(_03179_),
    .A2(_02814_),
    .A3(_02815_),
    .A4(_03101_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08397_ (.A1(_03102_),
    .A2(_03349_),
    .B(_01189_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08398_ (.A1(_01842_),
    .A2(_03348_),
    .A3(_03287_),
    .B(_03350_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08399_ (.A1(_03289_),
    .A2(_03346_),
    .B1(_03351_),
    .B2(_03055_),
    .C(_03211_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08400_ (.I(_02797_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08401_ (.I(_01892_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08402_ (.A1(_01841_),
    .A2(_01031_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08403_ (.A1(_03353_),
    .A2(_03354_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08404_ (.A1(_02800_),
    .A2(_01893_),
    .A3(_01032_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08405_ (.A1(_03355_),
    .A2(_03356_),
    .B(_01133_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08406_ (.I(_03334_),
    .Z(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08407_ (.A1(_03358_),
    .A2(_01895_),
    .B(_01161_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08408_ (.I(_03174_),
    .Z(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08409_ (.I(_03360_),
    .Z(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08410_ (.I(_03135_),
    .Z(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08411_ (.I(_03141_),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08412_ (.I(_03228_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08413_ (.I(_03232_),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08414_ (.A1(\as2650.stack[4][1] ),
    .A2(_03364_),
    .B1(_03365_),
    .B2(\as2650.stack[5][1] ),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08415_ (.I(_03319_),
    .Z(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08416_ (.I(_03321_),
    .Z(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08417_ (.A1(\as2650.stack[7][1] ),
    .A2(_03367_),
    .B1(_03368_),
    .B2(\as2650.stack[6][1] ),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08418_ (.A1(_03363_),
    .A2(_03366_),
    .A3(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08419_ (.A1(\as2650.stack[0][1] ),
    .A2(_03324_),
    .B1(_03325_),
    .B2(\as2650.stack[1][1] ),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08420_ (.A1(\as2650.stack[3][1] ),
    .A2(_03367_),
    .B1(_03368_),
    .B2(\as2650.stack[2][1] ),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08421_ (.A1(_03313_),
    .A2(_03371_),
    .A3(_03372_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08422_ (.A1(_03370_),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08423_ (.A1(\as2650.stack[11][1] ),
    .A2(_03220_),
    .B1(_03223_),
    .B2(\as2650.stack[10][1] ),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08424_ (.A1(\as2650.stack[8][1] ),
    .A2(_03229_),
    .B1(_03233_),
    .B2(\as2650.stack[9][1] ),
    .C(_03141_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08425_ (.A1(\as2650.stack[15][1] ),
    .A2(_03220_),
    .B1(_03223_),
    .B2(\as2650.stack[14][1] ),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08426_ (.A1(\as2650.stack[12][1] ),
    .A2(_03229_),
    .B1(_03233_),
    .B2(\as2650.stack[13][1] ),
    .C(_03246_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08427_ (.A1(_03375_),
    .A2(_03376_),
    .B1(_03377_),
    .B2(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08428_ (.A1(_03136_),
    .A2(_03379_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08429_ (.A1(_03362_),
    .A2(_03374_),
    .B(_03380_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08430_ (.A1(_03361_),
    .A2(_03381_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08431_ (.A1(_01895_),
    .A2(_03176_),
    .B(_03382_),
    .C(_03338_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08432_ (.A1(_03357_),
    .A2(_03359_),
    .B(_03256_),
    .C(_03383_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08433_ (.A1(_03353_),
    .A2(_03171_),
    .B(_03384_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08434_ (.A1(_02838_),
    .A2(_03295_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08435_ (.A1(_03299_),
    .A2(_01895_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08436_ (.A1(_03348_),
    .A2(_03385_),
    .B(_03387_),
    .C(_03193_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08437_ (.A1(_03386_),
    .A2(_03388_),
    .B(_03187_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08438_ (.A1(_03352_),
    .A2(_03385_),
    .B(_03389_),
    .C(_03289_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08439_ (.A1(_01046_),
    .A2(_03287_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08440_ (.I(_03391_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08441_ (.A1(_02846_),
    .A2(_03103_),
    .A3(_03102_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08442_ (.A1(_03387_),
    .A2(_03392_),
    .B1(_03393_),
    .B2(_03091_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08443_ (.A1(_03390_),
    .A2(_03394_),
    .B(_03028_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08444_ (.A1(_03098_),
    .A2(net91),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08445_ (.A1(_02862_),
    .A2(_03395_),
    .A3(_03106_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08446_ (.A1(_03287_),
    .A2(_03396_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08447_ (.I(_03089_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08448_ (.I(_03398_),
    .Z(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08449_ (.I(_03285_),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08450_ (.A1(_03400_),
    .A2(_01911_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08451_ (.A1(_03399_),
    .A2(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08452_ (.A1(_03067_),
    .A2(_03397_),
    .A3(_03402_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08453_ (.I(_01860_),
    .Z(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08454_ (.I(_03318_),
    .Z(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08455_ (.I(_03142_),
    .Z(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08456_ (.I(_03229_),
    .Z(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08457_ (.I(_03233_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08458_ (.A1(\as2650.stack[4][2] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\as2650.stack[5][2] ),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08459_ (.A1(\as2650.stack[7][2] ),
    .A2(_03221_),
    .B1(_03224_),
    .B2(\as2650.stack[6][2] ),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08460_ (.A1(_03406_),
    .A2(_03409_),
    .A3(_03410_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08461_ (.I(_03152_),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08462_ (.I(_03412_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08463_ (.A1(\as2650.stack[0][2] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\as2650.stack[1][2] ),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08464_ (.A1(\as2650.stack[3][2] ),
    .A2(_03221_),
    .B1(_03224_),
    .B2(\as2650.stack[2][2] ),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08465_ (.A1(_03413_),
    .A2(_03414_),
    .A3(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08466_ (.A1(_03411_),
    .A2(_03416_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08467_ (.I(_02589_),
    .Z(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08468_ (.I(_02671_),
    .Z(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08469_ (.A1(\as2650.stack[11][2] ),
    .A2(_03418_),
    .B1(_03419_),
    .B2(\as2650.stack[10][2] ),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08470_ (.I(_02634_),
    .Z(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08471_ (.A1(\as2650.stack[8][2] ),
    .A2(_03230_),
    .B1(_03421_),
    .B2(\as2650.stack[9][2] ),
    .C(_03363_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08472_ (.A1(\as2650.stack[15][2] ),
    .A2(_03418_),
    .B1(_03419_),
    .B2(\as2650.stack[14][2] ),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08473_ (.A1(\as2650.stack[12][2] ),
    .A2(_03230_),
    .B1(_03234_),
    .B2(\as2650.stack[13][2] ),
    .C(_03412_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08474_ (.A1(_03420_),
    .A2(_03422_),
    .B1(_03423_),
    .B2(_03424_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08475_ (.A1(_03305_),
    .A2(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08476_ (.A1(_03405_),
    .A2(_03417_),
    .B(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08477_ (.A1(_03360_),
    .A2(_03427_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08478_ (.I(_03302_),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08479_ (.A1(_01911_),
    .A2(_03429_),
    .B(_01160_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08480_ (.A1(_01132_),
    .A2(_01911_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08481_ (.A1(_01921_),
    .A2(_03355_),
    .Z(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08482_ (.A1(_03334_),
    .A2(_03432_),
    .B(_03337_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08483_ (.A1(_03428_),
    .A2(_03430_),
    .B1(_03431_),
    .B2(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08484_ (.A1(_03404_),
    .A2(_03434_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08485_ (.A1(_00571_),
    .A2(_03341_),
    .B(_03435_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08486_ (.A1(_00828_),
    .A2(_03397_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08487_ (.I(_03294_),
    .Z(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08488_ (.A1(_03347_),
    .A2(_03436_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08489_ (.A1(_03401_),
    .A2(_03439_),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08490_ (.I(_03294_),
    .Z(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08491_ (.A1(_02858_),
    .A2(_03441_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08492_ (.A1(_03438_),
    .A2(_03440_),
    .B(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08493_ (.A1(_01179_),
    .A2(_03437_),
    .B1(_03443_),
    .B2(_00512_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08494_ (.A1(_03352_),
    .A2(_03436_),
    .B1(_03444_),
    .B2(_01187_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08495_ (.A1(_03403_),
    .A2(_03445_),
    .B(_03028_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08496_ (.A1(_03108_),
    .A2(_03111_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08497_ (.A1(_03108_),
    .A2(_03111_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08498_ (.A1(_03182_),
    .A2(_03447_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08499_ (.A1(\as2650.stack[4][3] ),
    .A2(_01880_),
    .B1(_02635_),
    .B2(\as2650.stack[5][3] ),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08500_ (.I(_03319_),
    .Z(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08501_ (.I(_03321_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08502_ (.A1(\as2650.stack[7][3] ),
    .A2(_03450_),
    .B1(_03451_),
    .B2(\as2650.stack[6][3] ),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08503_ (.A1(_03363_),
    .A2(_03449_),
    .A3(_03452_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08504_ (.I(_01879_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08505_ (.A1(\as2650.stack[0][3] ),
    .A2(_03454_),
    .B1(_02635_),
    .B2(\as2650.stack[1][3] ),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08506_ (.A1(\as2650.stack[3][3] ),
    .A2(_03450_),
    .B1(_03451_),
    .B2(\as2650.stack[2][3] ),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08507_ (.A1(_03313_),
    .A2(_03455_),
    .A3(_03456_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08508_ (.A1(_03453_),
    .A2(_03457_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08509_ (.I(_03319_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08510_ (.I(_03321_),
    .Z(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08511_ (.A1(\as2650.stack[11][3] ),
    .A2(_03459_),
    .B1(_03460_),
    .B2(\as2650.stack[10][3] ),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08512_ (.I(_03228_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08513_ (.I(_03232_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08514_ (.A1(\as2650.stack[8][3] ),
    .A2(_03462_),
    .B1(_03463_),
    .B2(\as2650.stack[9][3] ),
    .C(_03241_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08515_ (.A1(\as2650.stack[15][3] ),
    .A2(_03367_),
    .B1(_03368_),
    .B2(\as2650.stack[14][3] ),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08516_ (.A1(\as2650.stack[12][3] ),
    .A2(_03462_),
    .B1(_03463_),
    .B2(\as2650.stack[13][3] ),
    .C(_03153_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08517_ (.A1(_03461_),
    .A2(_03464_),
    .B1(_03465_),
    .B2(_03466_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08518_ (.A1(_03318_),
    .A2(_03467_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08519_ (.A1(_03305_),
    .A2(_03458_),
    .B(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08520_ (.A1(_03360_),
    .A2(_03469_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08521_ (.A1(_01925_),
    .A2(_03429_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08522_ (.A1(_03337_),
    .A2(_03470_),
    .A3(_03471_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08523_ (.I(_01130_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08524_ (.A1(_01921_),
    .A2(\as2650.PC[3] ),
    .A3(_03355_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08525_ (.A1(_01921_),
    .A2(_03355_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08526_ (.A1(_01920_),
    .A2(_03475_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08527_ (.A1(_03474_),
    .A2(_03476_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08528_ (.A1(_01131_),
    .A2(_01924_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08529_ (.A1(_03473_),
    .A2(_03477_),
    .B(_03478_),
    .C(_01160_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08530_ (.A1(_03169_),
    .A2(_03472_),
    .A3(_03479_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08531_ (.A1(_01920_),
    .A2(_03170_),
    .B(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08532_ (.A1(_03285_),
    .A2(_01925_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08533_ (.A1(_03298_),
    .A2(_03481_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08534_ (.A1(_03294_),
    .A2(_03482_),
    .A3(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08535_ (.A1(_02873_),
    .A2(_03300_),
    .B(_03484_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08536_ (.A1(_02797_),
    .A2(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08537_ (.A1(_03296_),
    .A2(_03481_),
    .B(_03486_),
    .C(_03288_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08538_ (.A1(_03291_),
    .A2(_01925_),
    .A3(_03391_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08539_ (.A1(_03446_),
    .A2(_03448_),
    .B(_03487_),
    .C(_03488_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08540_ (.A1(_01308_),
    .A2(_03489_),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08541_ (.I(_03490_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08542_ (.A1(_03114_),
    .A2(_03099_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08543_ (.A1(_03113_),
    .A2(_03491_),
    .B(_03089_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08544_ (.A1(_03113_),
    .A2(_03491_),
    .B(_03492_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08545_ (.A1(_03286_),
    .A2(_01942_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08546_ (.A1(_03399_),
    .A2(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08547_ (.A1(_03049_),
    .A2(_03493_),
    .A3(_03495_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08548_ (.A1(\as2650.stack[4][4] ),
    .A2(_03306_),
    .B1(_03307_),
    .B2(\as2650.stack[5][4] ),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08549_ (.A1(\as2650.stack[7][4] ),
    .A2(_02590_),
    .B1(_02672_),
    .B2(\as2650.stack[6][4] ),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08550_ (.A1(_03242_),
    .A2(_03497_),
    .A3(_03498_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08551_ (.A1(\as2650.stack[0][4] ),
    .A2(_03306_),
    .B1(_03307_),
    .B2(\as2650.stack[1][4] ),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08552_ (.A1(\as2650.stack[3][4] ),
    .A2(_03309_),
    .B1(_03310_),
    .B2(\as2650.stack[2][4] ),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08553_ (.A1(_03247_),
    .A2(_03500_),
    .A3(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08554_ (.A1(_03499_),
    .A2(_03502_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08555_ (.A1(\as2650.stack[11][4] ),
    .A2(_03320_),
    .B1(_03322_),
    .B2(\as2650.stack[10][4] ),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08556_ (.A1(\as2650.stack[8][4] ),
    .A2(_03364_),
    .B1(_03365_),
    .B2(\as2650.stack[9][4] ),
    .C(_03241_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08557_ (.A1(\as2650.stack[15][4] ),
    .A2(_03320_),
    .B1(_03322_),
    .B2(\as2650.stack[14][4] ),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08558_ (.A1(\as2650.stack[12][4] ),
    .A2(_03454_),
    .B1(_03365_),
    .B2(\as2650.stack[13][4] ),
    .C(_03153_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08559_ (.A1(_03504_),
    .A2(_03505_),
    .B1(_03506_),
    .B2(_03507_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08560_ (.A1(_03318_),
    .A2(_03508_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08561_ (.A1(_03137_),
    .A2(_03503_),
    .B(_03509_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08562_ (.A1(_03175_),
    .A2(_03510_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08563_ (.A1(_01942_),
    .A2(_03303_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08564_ (.A1(_01195_),
    .A2(_03511_),
    .A3(_03512_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08565_ (.A1(\as2650.PC[4] ),
    .A2(_03474_),
    .Z(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08566_ (.A1(_03473_),
    .A2(_01942_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08567_ (.A1(_01132_),
    .A2(_03514_),
    .B(_03515_),
    .C(_01160_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08568_ (.A1(_03170_),
    .A2(_03513_),
    .A3(_03516_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08569_ (.A1(_01938_),
    .A2(_03256_),
    .B(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08570_ (.A1(_00828_),
    .A2(_03493_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08571_ (.A1(_03347_),
    .A2(_03518_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08572_ (.A1(_03441_),
    .A2(_03494_),
    .A3(_03520_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08573_ (.A1(_02887_),
    .A2(_03189_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08574_ (.A1(_03521_),
    .A2(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08575_ (.A1(_01179_),
    .A2(_03519_),
    .B1(_03523_),
    .B2(_00512_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08576_ (.A1(_03352_),
    .A2(_03518_),
    .B1(_03524_),
    .B2(_01187_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08577_ (.I(_02820_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08578_ (.A1(_03496_),
    .A2(_03525_),
    .B(_03526_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08579_ (.I(_02797_),
    .Z(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08580_ (.I(_03404_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08581_ (.I(_03362_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08582_ (.I(_02635_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08583_ (.A1(\as2650.stack[4][5] ),
    .A2(_01881_),
    .B1(_03530_),
    .B2(\as2650.stack[5][5] ),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08584_ (.I(_03450_),
    .Z(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08585_ (.I(_03451_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08586_ (.A1(\as2650.stack[7][5] ),
    .A2(_03532_),
    .B1(_03533_),
    .B2(\as2650.stack[6][5] ),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08587_ (.A1(_03243_),
    .A2(_03531_),
    .A3(_03534_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08588_ (.A1(\as2650.stack[0][5] ),
    .A2(_01881_),
    .B1(_02636_),
    .B2(\as2650.stack[1][5] ),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08589_ (.I(_03450_),
    .Z(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08590_ (.I(_03451_),
    .Z(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08591_ (.A1(\as2650.stack[3][5] ),
    .A2(_03537_),
    .B1(_03538_),
    .B2(\as2650.stack[2][5] ),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08592_ (.A1(_03413_),
    .A2(_03536_),
    .A3(_03539_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08593_ (.A1(_03535_),
    .A2(_03540_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08594_ (.I(_03459_),
    .Z(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08595_ (.I(_03460_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08596_ (.A1(\as2650.stack[11][5] ),
    .A2(_03542_),
    .B1(_03543_),
    .B2(\as2650.stack[10][5] ),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08597_ (.I(_03324_),
    .Z(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08598_ (.I(_03325_),
    .Z(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08599_ (.A1(\as2650.stack[8][5] ),
    .A2(_03545_),
    .B1(_03546_),
    .B2(\as2650.stack[9][5] ),
    .C(_03242_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08600_ (.A1(\as2650.stack[15][5] ),
    .A2(_03221_),
    .B1(_03224_),
    .B2(\as2650.stack[14][5] ),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08601_ (.A1(\as2650.stack[12][5] ),
    .A2(_03545_),
    .B1(_03546_),
    .B2(\as2650.stack[13][5] ),
    .C(_03247_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08602_ (.A1(_03544_),
    .A2(_03547_),
    .B1(_03548_),
    .B2(_03549_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08603_ (.A1(_03405_),
    .A2(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08604_ (.A1(_03529_),
    .A2(_03541_),
    .B(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08605_ (.A1(_03361_),
    .A2(_03552_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08606_ (.I(_03429_),
    .Z(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08607_ (.I(_01159_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08608_ (.A1(_01958_),
    .A2(_03554_),
    .B(_03555_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08609_ (.I(_01131_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08610_ (.A1(_03557_),
    .A2(_01958_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08611_ (.A1(_01938_),
    .A2(_03474_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08612_ (.A1(_01955_),
    .A2(_03559_),
    .Z(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08613_ (.A1(_03335_),
    .A2(_03560_),
    .B(_01195_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08614_ (.A1(_03553_),
    .A2(_03556_),
    .B1(_03558_),
    .B2(_03561_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08615_ (.A1(_03528_),
    .A2(_03562_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08616_ (.A1(_00560_),
    .A2(_03342_),
    .B(_03563_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08617_ (.A1(_02917_),
    .A2(_03295_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08618_ (.I(_03298_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08619_ (.A1(_03286_),
    .A2(_01958_),
    .Z(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08620_ (.A1(_03566_),
    .A2(_03564_),
    .B(_03567_),
    .C(_03193_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08621_ (.A1(_03565_),
    .A2(_03568_),
    .B(_03217_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08622_ (.I(_03288_),
    .Z(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08623_ (.A1(_03527_),
    .A2(_03564_),
    .B(_03569_),
    .C(_03570_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08624_ (.A1(_03116_),
    .A2(_03120_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08625_ (.I(_03398_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08626_ (.A1(_03116_),
    .A2(_03120_),
    .B(_01046_),
    .C(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08627_ (.A1(_03392_),
    .A2(_03567_),
    .B1(_03572_),
    .B2(_03574_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08628_ (.A1(_03571_),
    .A2(_03575_),
    .B(_03526_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08629_ (.A1(\as2650.stack[4][6] ),
    .A2(_03230_),
    .B1(_03234_),
    .B2(\as2650.stack[5][6] ),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08630_ (.I(_02589_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08631_ (.I(_02671_),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08632_ (.A1(\as2650.stack[7][6] ),
    .A2(_03577_),
    .B1(_03578_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08633_ (.A1(_03406_),
    .A2(_03576_),
    .A3(_03579_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08634_ (.I(_01879_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08635_ (.A1(\as2650.stack[0][6] ),
    .A2(_03581_),
    .B1(_03234_),
    .B2(\as2650.stack[1][6] ),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08636_ (.A1(\as2650.stack[3][6] ),
    .A2(_03577_),
    .B1(_03578_),
    .B2(\as2650.stack[2][6] ),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08637_ (.A1(_03154_),
    .A2(_03582_),
    .A3(_03583_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08638_ (.A1(_03580_),
    .A2(_03584_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08639_ (.A1(\as2650.stack[11][6] ),
    .A2(_02590_),
    .B1(_02672_),
    .B2(\as2650.stack[10][6] ),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08640_ (.I(_02634_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08641_ (.A1(\as2650.stack[8][6] ),
    .A2(_03454_),
    .B1(_03587_),
    .B2(\as2650.stack[9][6] ),
    .C(_03142_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08642_ (.A1(\as2650.stack[15][6] ),
    .A2(_03309_),
    .B1(_03310_),
    .B2(\as2650.stack[14][6] ),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08643_ (.A1(\as2650.stack[12][6] ),
    .A2(_01880_),
    .B1(_03587_),
    .B2(\as2650.stack[13][6] ),
    .C(_03412_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08644_ (.A1(_03586_),
    .A2(_03588_),
    .B1(_03589_),
    .B2(_03590_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08645_ (.A1(_03362_),
    .A2(_03591_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08646_ (.A1(_03137_),
    .A2(_03585_),
    .B(_03592_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08647_ (.A1(_01972_),
    .A2(_03304_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08648_ (.A1(_03304_),
    .A2(_03593_),
    .B(_03594_),
    .C(_01196_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08649_ (.A1(_01133_),
    .A2(_01972_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08650_ (.A1(_01938_),
    .A2(_00560_),
    .A3(_00557_),
    .A4(_03474_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08651_ (.A1(_01955_),
    .A2(_03559_),
    .B(_01969_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08652_ (.A1(_03597_),
    .A2(_03598_),
    .Z(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08653_ (.A1(_03358_),
    .A2(_03599_),
    .B(_03338_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08654_ (.A1(_03596_),
    .A2(_03600_),
    .B(_03039_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08655_ (.A1(_00557_),
    .A2(_03342_),
    .B1(_03595_),
    .B2(_03601_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08656_ (.A1(_02932_),
    .A2(_03295_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08657_ (.A1(_03299_),
    .A2(_01972_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08658_ (.A1(_03566_),
    .A2(_03602_),
    .B(_03604_),
    .C(_03189_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08659_ (.A1(_03603_),
    .A2(_03605_),
    .B(_03217_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08660_ (.A1(_03527_),
    .A2(_03602_),
    .B(_03606_),
    .C(_03570_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08661_ (.A1(_03097_),
    .A2(_03121_),
    .Z(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08662_ (.A1(_03392_),
    .A2(_03604_),
    .B1(_03608_),
    .B2(_03192_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08663_ (.A1(_03607_),
    .A2(_03609_),
    .B(_03526_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08664_ (.A1(_01981_),
    .A2(_03597_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08665_ (.A1(_01981_),
    .A2(_03597_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08666_ (.A1(_03557_),
    .A2(_03610_),
    .A3(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08667_ (.A1(_03358_),
    .A2(_01984_),
    .B(_03555_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08668_ (.A1(\as2650.stack[4][7] ),
    .A2(_03454_),
    .B1(_03587_),
    .B2(\as2650.stack[5][7] ),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08669_ (.A1(\as2650.stack[7][7] ),
    .A2(_03459_),
    .B1(_03460_),
    .B2(\as2650.stack[6][7] ),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08670_ (.A1(_03363_),
    .A2(_03614_),
    .A3(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08671_ (.A1(\as2650.stack[0][7] ),
    .A2(_03364_),
    .B1(_03587_),
    .B2(\as2650.stack[1][7] ),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08672_ (.A1(\as2650.stack[3][7] ),
    .A2(_03459_),
    .B1(_03460_),
    .B2(\as2650.stack[2][7] ),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08673_ (.A1(_03313_),
    .A2(_03617_),
    .A3(_03618_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08674_ (.A1(_03616_),
    .A2(_03619_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08675_ (.A1(\as2650.stack[11][7] ),
    .A2(_03367_),
    .B1(_03368_),
    .B2(\as2650.stack[10][7] ),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08676_ (.A1(\as2650.stack[8][7] ),
    .A2(_03462_),
    .B1(_03463_),
    .B2(\as2650.stack[9][7] ),
    .C(_03141_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08677_ (.A1(\as2650.stack[15][7] ),
    .A2(_03220_),
    .B1(_03223_),
    .B2(\as2650.stack[14][7] ),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08678_ (.A1(\as2650.stack[12][7] ),
    .A2(_03462_),
    .B1(_03463_),
    .B2(\as2650.stack[13][7] ),
    .C(_03246_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08679_ (.A1(_03621_),
    .A2(_03622_),
    .B1(_03623_),
    .B2(_03624_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08680_ (.A1(_03136_),
    .A2(_03625_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08681_ (.A1(_03362_),
    .A2(_03620_),
    .B(_03626_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08682_ (.A1(_03175_),
    .A2(_03627_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08683_ (.A1(_01984_),
    .A2(_03176_),
    .B(_03628_),
    .C(_03338_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08684_ (.A1(_03612_),
    .A2(_03613_),
    .B(_03256_),
    .C(_03629_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08685_ (.A1(_01996_),
    .A2(_03171_),
    .B(_03630_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08686_ (.A1(_03438_),
    .A2(_02948_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08687_ (.A1(_03299_),
    .A2(_01984_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08688_ (.A1(_03566_),
    .A2(_03631_),
    .B(_03633_),
    .C(_03189_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08689_ (.A1(_03632_),
    .A2(_03634_),
    .B(_03217_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08690_ (.A1(_03527_),
    .A2(_03631_),
    .B(_03635_),
    .C(_03570_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08691_ (.A1(_02937_),
    .A2(_03096_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08692_ (.A1(_03637_),
    .A2(_03121_),
    .B(_03125_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _08693_ (.A1(_03123_),
    .A2(_03638_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08694_ (.A1(_03391_),
    .A2(_03633_),
    .B1(_03639_),
    .B2(_03192_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08695_ (.A1(_03636_),
    .A2(_03640_),
    .B(_03526_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08696_ (.A1(\as2650.stack[4][8] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\as2650.stack[5][8] ),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08697_ (.A1(\as2650.stack[7][8] ),
    .A2(_03418_),
    .B1(_03419_),
    .B2(\as2650.stack[6][8] ),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08698_ (.A1(_03406_),
    .A2(_03641_),
    .A3(_03642_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08699_ (.A1(\as2650.stack[0][8] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\as2650.stack[1][8] ),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08700_ (.A1(\as2650.stack[3][8] ),
    .A2(_03418_),
    .B1(_03419_),
    .B2(\as2650.stack[2][8] ),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08701_ (.A1(_03413_),
    .A2(_03644_),
    .A3(_03645_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08702_ (.A1(_03643_),
    .A2(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08703_ (.A1(\as2650.stack[11][8] ),
    .A2(_03577_),
    .B1(_03578_),
    .B2(\as2650.stack[10][8] ),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08704_ (.A1(\as2650.stack[8][8] ),
    .A2(_03581_),
    .B1(_03421_),
    .B2(\as2650.stack[9][8] ),
    .C(_03142_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08705_ (.A1(\as2650.stack[15][8] ),
    .A2(_03577_),
    .B1(_03578_),
    .B2(\as2650.stack[14][8] ),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08706_ (.A1(\as2650.stack[12][8] ),
    .A2(_03581_),
    .B1(_03421_),
    .B2(\as2650.stack[13][8] ),
    .C(_03412_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08707_ (.A1(_03648_),
    .A2(_03649_),
    .B1(_03650_),
    .B2(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08708_ (.A1(_03305_),
    .A2(_03652_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08709_ (.A1(_03405_),
    .A2(_03647_),
    .B(_03653_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08710_ (.A1(_03360_),
    .A2(_03654_),
    .Z(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08711_ (.I(_01159_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08712_ (.A1(_01999_),
    .A2(_03303_),
    .B(_03655_),
    .C(_03656_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08713_ (.A1(_02000_),
    .A2(_03610_),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08714_ (.A1(_02000_),
    .A2(_03610_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08715_ (.A1(_03473_),
    .A2(_03659_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08716_ (.A1(_01132_),
    .A2(_01999_),
    .B1(_03658_),
    .B2(_03660_),
    .C(_03337_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08717_ (.A1(_02000_),
    .A2(_03404_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08718_ (.A1(_03404_),
    .A2(_03657_),
    .A3(_03661_),
    .B(_03662_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08719_ (.A1(_03347_),
    .A2(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08720_ (.A1(_03400_),
    .A2(_01999_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08721_ (.A1(_03300_),
    .A2(_03664_),
    .A3(_03665_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08722_ (.A1(_02971_),
    .A2(_03438_),
    .B(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08723_ (.A1(_03092_),
    .A2(_03128_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08724_ (.A1(_03398_),
    .A2(_03668_),
    .B(_00828_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08725_ (.A1(_00512_),
    .A2(_03667_),
    .B1(_03669_),
    .B2(_01179_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08726_ (.A1(_03352_),
    .A2(_03663_),
    .B1(_03670_),
    .B2(_01305_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08727_ (.A1(_03573_),
    .A2(_03665_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08728_ (.A1(_03399_),
    .A2(_03668_),
    .B(_03672_),
    .C(_03049_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08729_ (.I(_02820_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08730_ (.A1(_03671_),
    .A2(_03673_),
    .B(_03674_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08731_ (.A1(_03092_),
    .A2(_03128_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08732_ (.A1(_02977_),
    .A2(_03675_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08733_ (.A1(_03298_),
    .A2(_02013_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08734_ (.A1(_03573_),
    .A2(_03677_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08735_ (.A1(_03399_),
    .A2(_03676_),
    .B(_03678_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08736_ (.A1(_03341_),
    .A2(_03660_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08737_ (.A1(_02013_),
    .A2(_03554_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08738_ (.I(_03137_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08739_ (.I(_03581_),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08740_ (.I(_03421_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08741_ (.A1(\as2650.stack[4][9] ),
    .A2(_03683_),
    .B1(_03684_),
    .B2(\as2650.stack[5][9] ),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08742_ (.I(_02590_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08743_ (.A1(\as2650.stack[7][9] ),
    .A2(_03686_),
    .B1(_02673_),
    .B2(\as2650.stack[6][9] ),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08744_ (.A1(_03144_),
    .A2(_03685_),
    .A3(_03687_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08745_ (.A1(\as2650.stack[0][9] ),
    .A2(_03683_),
    .B1(_03684_),
    .B2(\as2650.stack[1][9] ),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08746_ (.I(_02672_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08747_ (.A1(\as2650.stack[3][9] ),
    .A2(_03686_),
    .B1(_03690_),
    .B2(\as2650.stack[2][9] ),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08748_ (.A1(_03248_),
    .A2(_03689_),
    .A3(_03691_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08749_ (.A1(_03688_),
    .A2(_03692_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08750_ (.A1(\as2650.stack[11][9] ),
    .A2(_03537_),
    .B1(_03538_),
    .B2(\as2650.stack[10][9] ),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08751_ (.I(_03364_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08752_ (.I(_03365_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08753_ (.A1(\as2650.stack[8][9] ),
    .A2(_03695_),
    .B1(_03696_),
    .B2(\as2650.stack[9][9] ),
    .C(_03143_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08754_ (.A1(\as2650.stack[15][9] ),
    .A2(_03537_),
    .B1(_03538_),
    .B2(\as2650.stack[14][9] ),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08755_ (.A1(\as2650.stack[12][9] ),
    .A2(_03695_),
    .B1(_03696_),
    .B2(\as2650.stack[13][9] ),
    .C(_03154_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08756_ (.A1(_03694_),
    .A2(_03697_),
    .B1(_03698_),
    .B2(_03699_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08757_ (.A1(_03529_),
    .A2(_03700_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08758_ (.A1(_03682_),
    .A2(_03693_),
    .B(_03701_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08759_ (.A1(_03361_),
    .A2(_03702_),
    .B(_03656_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08760_ (.A1(_03557_),
    .A2(_02013_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08761_ (.A1(_02014_),
    .A2(_03659_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08762_ (.A1(_03335_),
    .A2(_03705_),
    .B(_01195_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08763_ (.A1(_03681_),
    .A2(_03703_),
    .B1(_03704_),
    .B2(_03706_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08764_ (.A1(_02014_),
    .A2(_03680_),
    .B1(_03707_),
    .B2(_03528_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08765_ (.A1(_02807_),
    .A2(_03300_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08766_ (.A1(_03566_),
    .A2(_03708_),
    .B(_03677_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08767_ (.A1(_02982_),
    .A2(_03709_),
    .B1(_03710_),
    .B2(_03438_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08768_ (.I0(_03708_),
    .I1(_03711_),
    .S(_03073_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08769_ (.A1(_03055_),
    .A2(_03679_),
    .B1(_03712_),
    .B2(_03289_),
    .C(_03211_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08770_ (.A1(\as2650.stack[4][10] ),
    .A2(_03231_),
    .B1(_03235_),
    .B2(\as2650.stack[5][10] ),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08771_ (.A1(\as2650.stack[7][10] ),
    .A2(_02591_),
    .B1(_02673_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08772_ (.A1(_03144_),
    .A2(_03713_),
    .A3(_03714_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08773_ (.A1(\as2650.stack[0][10] ),
    .A2(_03683_),
    .B1(_03684_),
    .B2(\as2650.stack[1][10] ),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08774_ (.A1(\as2650.stack[3][10] ),
    .A2(_02591_),
    .B1(_02673_),
    .B2(\as2650.stack[2][10] ),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08775_ (.A1(_03155_),
    .A2(_03716_),
    .A3(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08776_ (.A1(_03715_),
    .A2(_03718_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08777_ (.A1(\as2650.stack[11][10] ),
    .A2(_02591_),
    .B1(_03690_),
    .B2(\as2650.stack[10][10] ),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08778_ (.A1(\as2650.stack[8][10] ),
    .A2(_01881_),
    .B1(_02636_),
    .B2(\as2650.stack[9][10] ),
    .C(_03406_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08779_ (.A1(\as2650.stack[15][10] ),
    .A2(_03686_),
    .B1(_03690_),
    .B2(\as2650.stack[14][10] ),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08780_ (.I(_03306_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08781_ (.A1(\as2650.stack[12][10] ),
    .A2(_03723_),
    .B1(_02636_),
    .B2(\as2650.stack[13][10] ),
    .C(_03413_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08782_ (.A1(_03720_),
    .A2(_03721_),
    .B1(_03722_),
    .B2(_03724_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08783_ (.A1(_03529_),
    .A2(_03725_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08784_ (.A1(_03682_),
    .A2(_03719_),
    .B(_03726_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08785_ (.I0(_02028_),
    .I1(_03727_),
    .S(_03175_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08786_ (.A1(_02014_),
    .A2(\as2650.PC[10] ),
    .A3(_03659_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08787_ (.A1(_02024_),
    .A2(_03705_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08788_ (.A1(_03729_),
    .A2(_03730_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08789_ (.A1(_03334_),
    .A2(_02027_),
    .B(_03656_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08790_ (.A1(_03335_),
    .A2(_03731_),
    .B(_03732_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08791_ (.A1(_01196_),
    .A2(_03728_),
    .B(_03733_),
    .C(_03039_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08792_ (.A1(_02024_),
    .A2(_03342_),
    .B(_03734_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08793_ (.A1(_03400_),
    .A2(_02028_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08794_ (.I(_03736_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08795_ (.A1(_03348_),
    .A2(_03735_),
    .B(_03737_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08796_ (.A1(_03190_),
    .A2(_03738_),
    .B(_03296_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08797_ (.A1(_02923_),
    .A2(_03193_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08798_ (.A1(_02996_),
    .A2(_03740_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08799_ (.A1(_03187_),
    .A2(_03735_),
    .B1(_03739_),
    .B2(_03741_),
    .C(_03288_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08800_ (.A1(_03092_),
    .A2(_02977_),
    .A3(_03128_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08801_ (.A1(_02850_),
    .A2(_03743_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08802_ (.A1(_03192_),
    .A2(_03744_),
    .B1(_03737_),
    .B2(_03392_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08803_ (.A1(_03742_),
    .A2(_03745_),
    .B(_03674_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08804_ (.A1(_02999_),
    .A2(_03129_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08805_ (.A1(_03091_),
    .A2(_03746_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08806_ (.A1(_03400_),
    .A2(_02041_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08807_ (.I(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08808_ (.I(_01532_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08809_ (.A1(_03358_),
    .A2(_03729_),
    .B(_03341_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08810_ (.A1(_02040_),
    .A2(_03554_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08811_ (.A1(\as2650.stack[4][11] ),
    .A2(_03683_),
    .B1(_03684_),
    .B2(\as2650.stack[5][11] ),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08812_ (.A1(\as2650.stack[7][11] ),
    .A2(_03686_),
    .B1(_03690_),
    .B2(\as2650.stack[6][11] ),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08813_ (.A1(_03243_),
    .A2(_03753_),
    .A3(_03754_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08814_ (.A1(\as2650.stack[0][11] ),
    .A2(_03723_),
    .B1(_03530_),
    .B2(\as2650.stack[1][11] ),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08815_ (.A1(\as2650.stack[3][11] ),
    .A2(_03532_),
    .B1(_03533_),
    .B2(\as2650.stack[2][11] ),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08816_ (.A1(_03248_),
    .A2(_03756_),
    .A3(_03757_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08817_ (.A1(_03755_),
    .A2(_03758_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08818_ (.A1(\as2650.stack[11][11] ),
    .A2(_03537_),
    .B1(_03538_),
    .B2(\as2650.stack[10][11] ),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08819_ (.A1(\as2650.stack[8][11] ),
    .A2(_03695_),
    .B1(_03696_),
    .B2(\as2650.stack[9][11] ),
    .C(_03143_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08820_ (.A1(\as2650.stack[15][11] ),
    .A2(_03542_),
    .B1(_03543_),
    .B2(\as2650.stack[14][11] ),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08821_ (.A1(\as2650.stack[12][11] ),
    .A2(_03695_),
    .B1(_03696_),
    .B2(\as2650.stack[13][11] ),
    .C(_03154_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08822_ (.A1(_03760_),
    .A2(_03761_),
    .B1(_03762_),
    .B2(_03763_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08823_ (.A1(_03529_),
    .A2(_03764_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08824_ (.A1(_03682_),
    .A2(_03759_),
    .B(_03765_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08825_ (.A1(_03361_),
    .A2(_03766_),
    .B(_03656_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08826_ (.A1(_02038_),
    .A2(_03729_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08827_ (.A1(_01131_),
    .A2(_03768_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08828_ (.A1(_03557_),
    .A2(_02040_),
    .B(_03769_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08829_ (.A1(_03752_),
    .A2(_03767_),
    .B1(_03770_),
    .B2(_03555_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08830_ (.A1(_02037_),
    .A2(_03751_),
    .B1(_03771_),
    .B2(_03039_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08831_ (.A1(_03291_),
    .A2(_03772_),
    .B(_03748_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08832_ (.A1(_03003_),
    .A2(_03709_),
    .B1(_03773_),
    .B2(_03441_),
    .C(_01532_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08833_ (.A1(_03750_),
    .A2(_03772_),
    .B(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08834_ (.A1(_03391_),
    .A2(_03749_),
    .B1(_03775_),
    .B2(_03289_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08835_ (.A1(_03747_),
    .A2(_03776_),
    .B(_03674_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08836_ (.A1(_03473_),
    .A2(_02050_),
    .B(_03769_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08837_ (.A1(_02052_),
    .A2(_03777_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08838_ (.A1(_02052_),
    .A2(_02050_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08839_ (.A1(\as2650.stack[4][12] ),
    .A2(_03723_),
    .B1(_03530_),
    .B2(\as2650.stack[5][12] ),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08840_ (.A1(\as2650.stack[7][12] ),
    .A2(_03532_),
    .B1(_03533_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08841_ (.A1(_03243_),
    .A2(_03780_),
    .A3(_03781_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08842_ (.A1(\as2650.stack[0][12] ),
    .A2(_03723_),
    .B1(_03530_),
    .B2(\as2650.stack[1][12] ),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08843_ (.A1(\as2650.stack[3][12] ),
    .A2(_03532_),
    .B1(_03533_),
    .B2(\as2650.stack[2][12] ),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08844_ (.A1(_03248_),
    .A2(_03783_),
    .A3(_03784_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08845_ (.A1(_03782_),
    .A2(_03785_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08846_ (.A1(\as2650.stack[11][12] ),
    .A2(_03542_),
    .B1(_03543_),
    .B2(\as2650.stack[10][12] ),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08847_ (.A1(\as2650.stack[8][12] ),
    .A2(_03545_),
    .B1(_03546_),
    .B2(\as2650.stack[9][12] ),
    .C(_03143_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08848_ (.A1(\as2650.stack[15][12] ),
    .A2(_03542_),
    .B1(_03543_),
    .B2(\as2650.stack[14][12] ),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08849_ (.A1(\as2650.stack[12][12] ),
    .A2(_03545_),
    .B1(_03546_),
    .B2(\as2650.stack[13][12] ),
    .C(_03247_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08850_ (.A1(_03787_),
    .A2(_03788_),
    .B1(_03789_),
    .B2(_03790_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08851_ (.A1(_03405_),
    .A2(_03791_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08852_ (.A1(_03682_),
    .A2(_03786_),
    .B(_03792_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08853_ (.A1(_03303_),
    .A2(_03793_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08854_ (.A1(_03779_),
    .A2(_03554_),
    .B(_03794_),
    .C(_03555_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08855_ (.A1(_01161_),
    .A2(_03778_),
    .B(_03795_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08856_ (.A1(_02052_),
    .A2(_03528_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08857_ (.A1(_03528_),
    .A2(_03796_),
    .B(_03797_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08858_ (.A1(_03286_),
    .A2(_03779_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08859_ (.A1(_03291_),
    .A2(_03798_),
    .B(_03799_),
    .C(_03441_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08860_ (.A1(_03012_),
    .A2(_03740_),
    .B(_03800_),
    .C(_03296_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08861_ (.A1(_03527_),
    .A2(_03798_),
    .B(_03801_),
    .C(_03570_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08862_ (.A1(_02999_),
    .A2(_03129_),
    .B(_03007_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08863_ (.A1(_03398_),
    .A2(_02051_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08864_ (.A1(_03573_),
    .A2(_03130_),
    .A3(_03803_),
    .B1(_03804_),
    .B2(_03348_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08865_ (.A1(_03055_),
    .A2(_03805_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08866_ (.A1(_03802_),
    .A2(_03806_),
    .B(_03674_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08867_ (.I(_02521_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08868_ (.A1(_02524_),
    .A2(_02529_),
    .B(_03807_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08869_ (.I(_02518_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08870_ (.A1(_02516_),
    .A2(_03809_),
    .B(_02525_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08871_ (.A1(_01141_),
    .A2(_03810_),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08872_ (.A1(_01554_),
    .A2(_02110_),
    .B1(_02347_),
    .B2(_03808_),
    .C(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08873_ (.A1(_01156_),
    .A2(_02181_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08874_ (.I(_03813_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08875_ (.I(_03814_),
    .Z(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08876_ (.A1(_00660_),
    .A2(_01392_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08877_ (.A1(_01855_),
    .A2(_03816_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08878_ (.A1(_01151_),
    .A2(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08879_ (.A1(_01394_),
    .A2(_03818_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08880_ (.I(_02174_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08881_ (.I(_03820_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08882_ (.I(_00639_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08883_ (.I(_03822_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08884_ (.A1(_01135_),
    .A2(_02347_),
    .A3(_01210_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08885_ (.A1(_03823_),
    .A2(_03824_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08886_ (.A1(_03821_),
    .A2(_03825_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08887_ (.A1(_01146_),
    .A2(_02127_),
    .Z(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08888_ (.A1(_01391_),
    .A2(_03827_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08889_ (.I(_03828_),
    .Z(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08890_ (.A1(_03819_),
    .A2(_03826_),
    .A3(_03829_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08891_ (.I(_00666_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08892_ (.A1(_03831_),
    .A2(_01392_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08893_ (.A1(_01855_),
    .A2(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08894_ (.I(_01142_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08895_ (.A1(_03823_),
    .A2(_03821_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08896_ (.A1(_01143_),
    .A2(_02144_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08897_ (.A1(_03835_),
    .A2(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08898_ (.A1(_01068_),
    .A2(_01204_),
    .B(_01284_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08899_ (.A1(_03834_),
    .A2(_02153_),
    .A3(_03837_),
    .A4(_03838_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08900_ (.A1(_01857_),
    .A2(_03833_),
    .A3(_03839_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08901_ (.A1(_01194_),
    .A2(_01206_),
    .A3(_03169_),
    .A4(_03840_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08902_ (.A1(_02438_),
    .A2(_03815_),
    .B(_03830_),
    .C(_03841_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08903_ (.I(_03841_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08904_ (.I(_03843_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08905_ (.A1(_03831_),
    .A2(_01393_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08906_ (.A1(_01856_),
    .A2(_03845_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08907_ (.I(_03846_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08908_ (.A1(_01391_),
    .A2(_02130_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08909_ (.I(_02139_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08910_ (.I(_00795_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08911_ (.A1(_03850_),
    .A2(_02543_),
    .B(_01578_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(_01578_),
    .A2(_02152_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08913_ (.I(_02543_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08914_ (.A1(_02135_),
    .A2(_03851_),
    .B1(_03852_),
    .B2(_03853_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08915_ (.A1(_01555_),
    .A2(_03849_),
    .B(_03854_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08916_ (.A1(_03823_),
    .A2(_02186_),
    .A3(_03836_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08917_ (.I(_03856_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(_01554_),
    .A2(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08919_ (.A1(_01222_),
    .A2(_03857_),
    .B(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08920_ (.A1(_03853_),
    .A2(_02135_),
    .A3(_03859_),
    .B(_03848_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08921_ (.A1(_01147_),
    .A2(_03832_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08922_ (.A1(_03830_),
    .A2(_03861_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08923_ (.A1(_03848_),
    .A2(_03812_),
    .B1(_03855_),
    .B2(_03860_),
    .C(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08924_ (.A1(_03331_),
    .A2(_03847_),
    .B(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08925_ (.A1(_03844_),
    .A2(_03864_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08926_ (.A1(_01555_),
    .A2(_03842_),
    .B(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08927_ (.I(_03866_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08928_ (.A1(_01207_),
    .A2(_02172_),
    .A3(_03172_),
    .A4(_02354_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08929_ (.A1(_01289_),
    .A2(_03868_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08930_ (.A1(_02131_),
    .A2(_03869_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08931_ (.I(_03870_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08932_ (.A1(_01207_),
    .A2(_01208_),
    .A3(_01198_),
    .A4(_03172_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08933_ (.I(_03872_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08934_ (.I(_02130_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08935_ (.I(_03874_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08936_ (.A1(_03875_),
    .A2(_03812_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08937_ (.A1(_03875_),
    .A2(_03867_),
    .B(_03876_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08938_ (.I(_03821_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08939_ (.I(_03878_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08940_ (.A1(_03879_),
    .A2(_03867_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08941_ (.A1(_02177_),
    .A2(_03872_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08942_ (.I(_02187_),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08943_ (.I(_03882_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08944_ (.A1(_02089_),
    .A2(_01556_),
    .B(_03883_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08945_ (.A1(_03881_),
    .A2(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08946_ (.A1(_01555_),
    .A2(_02188_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08947_ (.I(_03823_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08948_ (.A1(_03887_),
    .A2(_03873_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08949_ (.A1(_02089_),
    .A2(_03886_),
    .B(_03888_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08950_ (.A1(_03885_),
    .A2(_03889_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08951_ (.A1(_03873_),
    .A2(_03877_),
    .B1(_03880_),
    .B2(_03890_),
    .C(_03870_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08952_ (.A1(_03867_),
    .A2(_03871_),
    .B(_03891_),
    .C(_02183_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08953_ (.I(_02939_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08954_ (.A1(_02183_),
    .A2(_03812_),
    .B(_03892_),
    .C(_03893_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08955_ (.A1(_01384_),
    .A2(_01114_),
    .A3(_01328_),
    .A4(_01137_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08956_ (.I(_03894_),
    .Z(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08957_ (.I(_03895_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08958_ (.I(_03878_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08959_ (.A1(_01288_),
    .A2(_03868_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08960_ (.A1(_03897_),
    .A2(_01176_),
    .A3(_03898_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08961_ (.A1(_01541_),
    .A2(_03896_),
    .A3(_03899_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _08962_ (.I(_01568_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08963_ (.A1(_03822_),
    .A2(_03836_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08964_ (.I(_03902_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08965_ (.A1(_03879_),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08966_ (.A1(_03861_),
    .A2(_03904_),
    .B(_03257_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08967_ (.I(_03847_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08968_ (.I(_03906_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08969_ (.I(_03857_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08970_ (.A1(_03381_),
    .A2(_03907_),
    .B1(_03908_),
    .B2(net84),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08971_ (.I(_03257_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08972_ (.A1(_03901_),
    .A2(_03905_),
    .B1(_03909_),
    .B2(_03910_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08973_ (.A1(_03900_),
    .A2(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08974_ (.I(_03887_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08975_ (.A1(_02228_),
    .A2(_03913_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08976_ (.A1(_02229_),
    .A2(_03901_),
    .B(_03900_),
    .C(_03914_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08977_ (.A1(_01184_),
    .A2(_03915_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08978_ (.A1(_03912_),
    .A2(_03916_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08979_ (.A1(_03807_),
    .A2(_02534_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08980_ (.A1(_02524_),
    .A2(_02535_),
    .B(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08981_ (.I(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08982_ (.I(_02110_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08983_ (.A1(_03029_),
    .A2(_03874_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08984_ (.A1(_03920_),
    .A2(_03921_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08985_ (.A1(_01914_),
    .A2(_03857_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08986_ (.A1(_01573_),
    .A2(_03908_),
    .B(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08987_ (.A1(_01139_),
    .A2(_03814_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08988_ (.A1(_03815_),
    .A2(_03924_),
    .B1(_03919_),
    .B2(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08989_ (.A1(_03427_),
    .A2(_03861_),
    .B1(_03862_),
    .B2(_03926_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08990_ (.A1(_03920_),
    .A2(_03815_),
    .B(_03830_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08991_ (.A1(_03844_),
    .A2(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08992_ (.A1(_01574_),
    .A2(_03929_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08993_ (.A1(_03841_),
    .A2(_03927_),
    .B(_03930_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08994_ (.A1(_03920_),
    .A2(_02182_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08995_ (.A1(_02301_),
    .A2(_01573_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08996_ (.A1(_02301_),
    .A2(_02177_),
    .B(_03933_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08997_ (.A1(_03897_),
    .A2(_03934_),
    .B(_03895_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08998_ (.A1(_03896_),
    .A2(_03932_),
    .B(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08999_ (.A1(_03870_),
    .A2(_03936_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09000_ (.A1(_03879_),
    .A2(_03935_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09001_ (.A1(_03918_),
    .A2(_03932_),
    .B(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09002_ (.A1(_03871_),
    .A2(_03939_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09003_ (.A1(_03931_),
    .A2(_03937_),
    .B(_03922_),
    .C(_03940_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09004_ (.A1(_03919_),
    .A2(_03922_),
    .B(_03941_),
    .C(_03893_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09005_ (.A1(_03469_),
    .A2(_03907_),
    .B1(_03908_),
    .B2(net99),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09006_ (.A1(_03849_),
    .A2(_03905_),
    .B1(_03942_),
    .B2(_03910_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09007_ (.A1(_03061_),
    .A2(_03913_),
    .B(_03873_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09008_ (.A1(_03062_),
    .A2(_03849_),
    .B(_03899_),
    .C(_03944_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09009_ (.A1(_03900_),
    .A2(_03943_),
    .B1(_03945_),
    .B2(_03750_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09010_ (.A1(_00510_),
    .A2(_03946_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09011_ (.I(_02213_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09012_ (.I(_03947_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09013_ (.A1(_03510_),
    .A2(_03907_),
    .B1(_03908_),
    .B2(net100),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09014_ (.A1(_03948_),
    .A2(_03905_),
    .B1(_03949_),
    .B2(_03910_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09015_ (.A1(_03064_),
    .A2(_03913_),
    .B(_03873_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09016_ (.A1(_03064_),
    .A2(_03948_),
    .B(_03899_),
    .C(_03951_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09017_ (.A1(_03900_),
    .A2(_03950_),
    .B1(_03952_),
    .B2(_03750_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09018_ (.A1(_00510_),
    .A2(_03953_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09019_ (.A1(_01324_),
    .A2(_02139_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09020_ (.A1(_03849_),
    .A2(_01504_),
    .B(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09021_ (.A1(_01073_),
    .A2(_01209_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09022_ (.A1(_01325_),
    .A2(_03856_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09023_ (.A1(net101),
    .A2(_03856_),
    .B(_03957_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09024_ (.A1(_01578_),
    .A2(_02420_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09025_ (.A1(_02135_),
    .A2(_03954_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09026_ (.A1(_03956_),
    .A2(_03958_),
    .B1(_03959_),
    .B2(_03960_),
    .C(_03853_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09027_ (.A1(_03853_),
    .A2(_03955_),
    .B(_03961_),
    .C(_03814_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09028_ (.A1(_02354_),
    .A2(_02400_),
    .A3(_02418_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09029_ (.A1(_03925_),
    .A2(_03963_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09030_ (.A1(_03962_),
    .A2(_03964_),
    .B(_03862_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09031_ (.A1(_03552_),
    .A2(_03906_),
    .B(_03965_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09032_ (.A1(_01325_),
    .A2(_03929_),
    .B1(_03966_),
    .B2(_03844_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(_02177_),
    .A2(_03894_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09034_ (.I0(_03967_),
    .I1(_03963_),
    .S(_03932_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09035_ (.A1(_03881_),
    .A2(_03969_),
    .B(_03869_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09036_ (.I(_03882_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09037_ (.A1(_02436_),
    .A2(_01592_),
    .B(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09038_ (.A1(_02915_),
    .A2(_01591_),
    .A3(_03971_),
    .A4(_03869_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09039_ (.A1(_03881_),
    .A2(_03972_),
    .B1(_03973_),
    .B2(_03888_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09040_ (.A1(_03879_),
    .A2(_03967_),
    .B(_03974_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09041_ (.A1(_01541_),
    .A2(_01177_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09042_ (.A1(_03968_),
    .A2(_03970_),
    .B(_03975_),
    .C(_03976_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09043_ (.A1(_03871_),
    .A2(_03967_),
    .B(_03977_),
    .C(_03922_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09044_ (.A1(_03920_),
    .A2(_03921_),
    .A3(_03963_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09045_ (.A1(_03211_),
    .A2(_03978_),
    .A3(_03979_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09046_ (.A1(_01061_),
    .A2(_01521_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09047_ (.A1(_02929_),
    .A2(_01513_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09048_ (.A1(_02300_),
    .A2(_01465_),
    .B1(_01476_),
    .B2(_03060_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09049_ (.A1(_02391_),
    .A2(_01485_),
    .B1(_01497_),
    .B2(_02434_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09050_ (.A1(_03981_),
    .A2(_03982_),
    .A3(_03983_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09051_ (.A1(_02435_),
    .A2(_01497_),
    .B1(_01513_),
    .B2(_02929_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09052_ (.A1(_03060_),
    .A2(_01476_),
    .B1(_01485_),
    .B2(_02391_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09053_ (.A1(_02299_),
    .A2(_01465_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09054_ (.A1(_02088_),
    .A2(_01425_),
    .B1(_01449_),
    .B2(_02227_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09055_ (.A1(_02088_),
    .A2(_01425_),
    .B1(_01449_),
    .B2(_02227_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09056_ (.I(_03989_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09057_ (.A1(_03986_),
    .A2(_03987_),
    .A3(_03988_),
    .A4(_03990_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09058_ (.A1(_03980_),
    .A2(_03984_),
    .A3(_03985_),
    .A4(_03991_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09059_ (.A1(_02180_),
    .A2(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09060_ (.I(_03985_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09061_ (.A1(_02227_),
    .A2(_01449_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09062_ (.A1(_03988_),
    .A2(_03995_),
    .B(_03987_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09063_ (.A1(_02300_),
    .A2(_01465_),
    .B1(_01476_),
    .B2(_02360_),
    .C(_03996_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09064_ (.A1(_03986_),
    .A2(_03997_),
    .B(_03983_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09065_ (.A1(_03994_),
    .A2(_03998_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09066_ (.A1(_03981_),
    .A2(_03999_),
    .B(_03980_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09067_ (.A1(_02513_),
    .A2(_01569_),
    .A3(_01521_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09068_ (.A1(_00529_),
    .A2(_01568_),
    .A3(_01521_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09069_ (.A1(_04000_),
    .A2(_04001_),
    .A3(_04002_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09070_ (.A1(_03841_),
    .A2(_03818_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09071_ (.A1(_03593_),
    .A2(_03847_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09072_ (.A1(_02486_),
    .A2(_02490_),
    .A3(_02492_),
    .B1(_02477_),
    .B2(_02303_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09073_ (.A1(_02125_),
    .A2(_02265_),
    .A3(_02325_),
    .A4(_02368_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09074_ (.A1(_02418_),
    .A2(_02457_),
    .A3(_04007_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09075_ (.A1(_04006_),
    .A2(_04008_),
    .B(_02534_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09076_ (.I(_02158_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09077_ (.A1(_00774_),
    .A2(_00765_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09078_ (.A1(_01079_),
    .A2(_04011_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09079_ (.A1(_03850_),
    .A2(_02142_),
    .A3(_02327_),
    .A4(_04012_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09080_ (.A1(_02146_),
    .A2(_02545_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09081_ (.A1(_01079_),
    .A2(_00848_),
    .A3(_02141_),
    .A4(_04011_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09082_ (.A1(_00779_),
    .A2(_03956_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09083_ (.A1(_03820_),
    .A2(_01272_),
    .B(_01122_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09084_ (.A1(_01083_),
    .A2(_03822_),
    .A3(_01119_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09085_ (.A1(_02144_),
    .A2(_04018_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09086_ (.A1(\as2650.debug_psu[4] ),
    .A2(\as2650.debug_psu[5] ),
    .A3(net144),
    .A4(_03132_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09087_ (.A1(_03820_),
    .A2(_04020_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09088_ (.A1(\as2650.debug_psl[6] ),
    .A2(_01349_),
    .A3(\as2650.debug_psl[0] ),
    .A4(\as2650.debug_psl[5] ),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09089_ (.A1(\as2650.debug_psl[1] ),
    .A2(\as2650.debug_psl[2] ),
    .A3(_01577_),
    .A4(_04022_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09090_ (.I(\as2650.debug_psl[7] ),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09091_ (.A1(_04024_),
    .A2(_01121_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09092_ (.A1(\as2650.debug_psu[7] ),
    .A2(_04021_),
    .B1(_04023_),
    .B2(_04025_),
    .C(_04019_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09093_ (.A1(_01319_),
    .A2(_04019_),
    .B(_04026_),
    .C(_03902_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09094_ (.A1(_03903_),
    .A2(_04017_),
    .B(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09095_ (.A1(_04015_),
    .A2(_04016_),
    .B1(_04028_),
    .B2(_03956_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09096_ (.A1(_04013_),
    .A2(_04014_),
    .B1(_04029_),
    .B2(_02146_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09097_ (.A1(_01259_),
    .A2(net101),
    .A3(_01273_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09098_ (.A1(net73),
    .A2(net84),
    .A3(net95),
    .A4(net99),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09099_ (.A1(_04031_),
    .A2(_04032_),
    .B(_01280_),
    .C(_04010_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09100_ (.A1(_04010_),
    .A2(_04030_),
    .B(_04033_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09101_ (.A1(_03813_),
    .A2(_04034_),
    .B(_03828_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09102_ (.A1(_03814_),
    .A2(_04009_),
    .B(_04035_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09103_ (.A1(_01060_),
    .A2(_01281_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09104_ (.A1(_03850_),
    .A2(_01987_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09105_ (.A1(_01503_),
    .A2(_01273_),
    .B(_04038_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _09106_ (.A1(_01096_),
    .A2(_01482_),
    .B1(_01961_),
    .B2(_01087_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09107_ (.A1(_01087_),
    .A2(_01961_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09108_ (.A1(_00893_),
    .A2(_01259_),
    .B(_04041_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09109_ (.A1(_01472_),
    .A2(_01928_),
    .B(_04040_),
    .C(_04042_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09110_ (.A1(_01456_),
    .A2(net95),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09111_ (.A1(_00847_),
    .A2(_01222_),
    .B1(_01442_),
    .B2(_01438_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09112_ (.A1(_01433_),
    .A2(_01236_),
    .B(_04045_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09113_ (.A1(_01456_),
    .A2(net95),
    .B1(_01251_),
    .B2(_01093_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09114_ (.A1(_04044_),
    .A2(_04046_),
    .B(_04047_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09115_ (.A1(_01503_),
    .A2(_01273_),
    .B1(_04040_),
    .B2(_04041_),
    .C1(_04043_),
    .C2(_04048_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09116_ (.A1(_01568_),
    .A2(_04038_),
    .B1(_04039_),
    .B2(_04049_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09117_ (.A1(_04037_),
    .A2(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09118_ (.A1(_03901_),
    .A2(_04037_),
    .B(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09119_ (.A1(_01101_),
    .A2(net73),
    .B1(net102),
    .B2(_01503_),
    .C1(net84),
    .C2(_01433_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09120_ (.A1(_01060_),
    .A2(_01280_),
    .B(_04039_),
    .C(_04044_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09121_ (.A1(_04047_),
    .A2(_04045_),
    .A3(_04053_),
    .A4(_04054_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09122_ (.A1(_04043_),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09123_ (.A1(_04052_),
    .A2(_04056_),
    .B(_03829_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09124_ (.A1(_04036_),
    .A2(_04057_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09125_ (.A1(_03887_),
    .A2(_02186_),
    .A3(_03824_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09126_ (.I(_01277_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09127_ (.A1(_04060_),
    .A2(_01338_),
    .B1(_01343_),
    .B2(_01258_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09128_ (.I(_04061_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09129_ (.A1(_01258_),
    .A2(_04060_),
    .A3(net75),
    .A4(_01344_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09130_ (.A1(_04062_),
    .A2(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09131_ (.A1(_01254_),
    .A2(_01330_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09132_ (.A1(_01239_),
    .A2(_01354_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09133_ (.A1(_04065_),
    .A2(_04066_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09134_ (.A1(_01262_),
    .A2(_01334_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09135_ (.A1(_04065_),
    .A2(_04066_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09136_ (.A1(_04067_),
    .A2(_04068_),
    .B(_04069_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09137_ (.I(_01331_),
    .Z(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09138_ (.I(_01354_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09139_ (.A1(_01248_),
    .A2(_01263_),
    .A3(_04071_),
    .A4(_04072_),
    .Z(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09140_ (.A1(_01263_),
    .A2(_01332_),
    .B1(_01355_),
    .B2(_01249_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09141_ (.A1(_04073_),
    .A2(_04074_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09142_ (.A1(_01269_),
    .A2(_01335_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09143_ (.A1(_04075_),
    .A2(_04076_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09144_ (.A1(_04070_),
    .A2(_04077_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09145_ (.A1(_04070_),
    .A2(_04077_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09146_ (.A1(_04078_),
    .A2(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09147_ (.A1(_04064_),
    .A2(_04080_),
    .B(_04078_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09148_ (.I(_04081_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09149_ (.A1(_01265_),
    .A2(_01344_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09150_ (.A1(_04075_),
    .A2(_04076_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09151_ (.A1(_04073_),
    .A2(_04084_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09152_ (.A1(_01253_),
    .A2(_01268_),
    .A3(_02067_),
    .A4(_02080_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09153_ (.A1(_01270_),
    .A2(net77),
    .B1(_01355_),
    .B2(_01257_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09154_ (.A1(_04086_),
    .A2(_04087_),
    .Z(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09155_ (.A1(_04060_),
    .A2(net76),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09156_ (.A1(_04088_),
    .A2(_04089_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09157_ (.A1(_04085_),
    .A2(_04090_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09158_ (.A1(_04083_),
    .A2(_04091_),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09159_ (.A1(_04082_),
    .A2(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09160_ (.A1(_04082_),
    .A2(_04092_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09161_ (.I(_04094_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09162_ (.A1(_04063_),
    .A2(_04095_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09163_ (.A1(_01271_),
    .A2(_01344_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09164_ (.A1(_01265_),
    .A2(_01278_),
    .A3(net77),
    .A4(net79),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09165_ (.A1(_01276_),
    .A2(_02067_),
    .B1(_02081_),
    .B2(_01961_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09166_ (.A1(_04098_),
    .A2(_04099_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09167_ (.A1(_04088_),
    .A2(_04089_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09168_ (.A1(_04086_),
    .A2(_04101_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09169_ (.A1(_04100_),
    .A2(_04102_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09170_ (.A1(_04097_),
    .A2(_04103_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09171_ (.A1(_01266_),
    .A2(net78),
    .A3(_04091_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09172_ (.A1(_04085_),
    .A2(_04090_),
    .B(_04105_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09173_ (.A1(_04104_),
    .A2(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09174_ (.A1(_04093_),
    .A2(_04096_),
    .B(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09175_ (.A1(_01279_),
    .A2(net78),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09176_ (.A1(_01268_),
    .A2(_02081_),
    .B(_04098_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09177_ (.A1(_01975_),
    .A2(_04098_),
    .B(_04110_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09178_ (.A1(_04109_),
    .A2(_04111_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09179_ (.A1(_01272_),
    .A2(net78),
    .A3(_04103_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09180_ (.A1(_04100_),
    .A2(_04102_),
    .B(_04113_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09181_ (.A1(_04112_),
    .A2(_04114_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09182_ (.A1(_04104_),
    .A2(_04106_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09183_ (.A1(_04116_),
    .A2(_04108_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09184_ (.A1(_04117_),
    .A2(_04115_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09185_ (.A1(_04063_),
    .A2(_04094_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09186_ (.A1(_01247_),
    .A2(_01330_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09187_ (.A1(_01231_),
    .A2(_01354_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09188_ (.A1(_04120_),
    .A2(_04121_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09189_ (.A1(_01255_),
    .A2(_01333_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09190_ (.A1(_04120_),
    .A2(_04121_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09191_ (.A1(_04122_),
    .A2(_04123_),
    .B(_04124_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09192_ (.A1(_04065_),
    .A2(_04066_),
    .A3(_04068_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09193_ (.A1(_04125_),
    .A2(_04126_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09194_ (.A1(_01246_),
    .A2(_02074_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09195_ (.I(_01336_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09196_ (.A1(_01269_),
    .A2(_04129_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09197_ (.I(_01340_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09198_ (.A1(_01277_),
    .A2(_04131_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09199_ (.A1(_04128_),
    .A2(_04130_),
    .A3(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09200_ (.I(_04126_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09201_ (.A1(_04125_),
    .A2(_04134_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09202_ (.A1(_04127_),
    .A2(_04133_),
    .B(_04135_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09203_ (.A1(_04064_),
    .A2(_04080_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09204_ (.A1(_04130_),
    .A2(_04132_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09205_ (.A1(_04130_),
    .A2(_04132_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09206_ (.A1(_04128_),
    .A2(_04138_),
    .B(_04139_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09207_ (.A1(_04136_),
    .A2(_04137_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09208_ (.A1(_04140_),
    .A2(_04141_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09209_ (.A1(_04136_),
    .A2(_04137_),
    .B(_04142_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09210_ (.A1(_04119_),
    .A2(_04143_),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09211_ (.A1(_01248_),
    .A2(_01334_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09212_ (.I(_01240_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09213_ (.A1(_04146_),
    .A2(_04071_),
    .B1(_04072_),
    .B2(_01224_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09214_ (.A1(_01225_),
    .A2(_04146_),
    .A3(_04071_),
    .A4(_04072_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09215_ (.A1(_04145_),
    .A2(_04147_),
    .B(_04148_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09216_ (.A1(_04120_),
    .A2(_04121_),
    .A3(_04123_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09217_ (.A1(_04149_),
    .A2(_04150_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09218_ (.A1(_01241_),
    .A2(_01343_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09219_ (.A1(_01269_),
    .A2(_01339_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09220_ (.A1(_01262_),
    .A2(_01336_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09221_ (.A1(_04153_),
    .A2(_04154_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09222_ (.A1(_04152_),
    .A2(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09223_ (.A1(_04149_),
    .A2(_04150_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09224_ (.A1(_04151_),
    .A2(_04156_),
    .B(_04157_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09225_ (.A1(_04127_),
    .A2(_04133_),
    .Z(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09226_ (.A1(_04158_),
    .A2(_04159_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09227_ (.A1(_01238_),
    .A2(_02074_),
    .A3(_04155_),
    .B1(_04154_),
    .B2(_04153_),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09228_ (.A1(_04158_),
    .A2(_04159_),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09229_ (.A1(_04161_),
    .A2(_04162_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09230_ (.A1(_04140_),
    .A2(_04141_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09231_ (.A1(_04160_),
    .A2(_04163_),
    .B(_04164_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09232_ (.A1(_04144_),
    .A2(_04165_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09233_ (.A1(_04164_),
    .A2(_04160_),
    .A3(_04163_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09234_ (.A1(_04165_),
    .A2(_04167_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09235_ (.I(_01340_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09236_ (.A1(_01256_),
    .A2(_01264_),
    .A3(_01337_),
    .A4(_04169_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09237_ (.A1(_01232_),
    .A2(_01343_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09238_ (.I(_04129_),
    .Z(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09239_ (.A1(_01256_),
    .A2(_04172_),
    .B1(_04169_),
    .B2(_01264_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09240_ (.A1(_04171_),
    .A2(_04170_),
    .A3(_04173_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09241_ (.A1(_04170_),
    .A2(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09242_ (.A1(_04060_),
    .A2(_01347_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09243_ (.A1(_04175_),
    .A2(_04176_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09244_ (.A1(_04175_),
    .A2(_04176_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09245_ (.A1(_04170_),
    .A2(_04173_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09246_ (.A1(_04171_),
    .A2(_04179_),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09247_ (.A1(_01231_),
    .A2(_01239_),
    .A3(_01330_),
    .A4(_01333_),
    .Z(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09248_ (.I(_04181_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09249_ (.A1(_01240_),
    .A2(_01331_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09250_ (.A1(_01224_),
    .A2(_04072_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09251_ (.A1(_04183_),
    .A2(_04184_),
    .A3(_04145_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09252_ (.A1(_04182_),
    .A2(_04185_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09253_ (.A1(_04182_),
    .A2(_04185_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09254_ (.A1(_04180_),
    .A2(_04186_),
    .B(_04187_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09255_ (.A1(_04151_),
    .A2(_04156_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09256_ (.A1(_04188_),
    .A2(_04189_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09257_ (.A1(_04188_),
    .A2(_04189_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09258_ (.A1(_04178_),
    .A2(_04190_),
    .B(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09259_ (.A1(_04161_),
    .A2(_04162_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09260_ (.A1(_04192_),
    .A2(_04193_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09261_ (.A1(_04192_),
    .A2(_04193_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09262_ (.A1(_04177_),
    .A2(_04194_),
    .B(_04195_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09263_ (.A1(_04168_),
    .A2(_04196_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09264_ (.A1(_01223_),
    .A2(_01342_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09265_ (.A1(_01249_),
    .A2(_01338_),
    .B1(_01341_),
    .B2(_01257_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09266_ (.A1(_01249_),
    .A2(_01257_),
    .A3(_04172_),
    .A4(_01341_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09267_ (.A1(_04198_),
    .A2(_04199_),
    .B(_04200_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09268_ (.A1(_01271_),
    .A2(net105),
    .A3(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09269_ (.A1(_01270_),
    .A2(_01346_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09270_ (.A1(_04201_),
    .A2(_04203_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09271_ (.A1(_01278_),
    .A2(_01353_),
    .A3(_04204_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09272_ (.A1(_04202_),
    .A2(_04205_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09273_ (.A1(_01278_),
    .A2(_01352_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09274_ (.A1(_04207_),
    .A2(_04204_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09275_ (.A1(_01233_),
    .A2(_04071_),
    .B1(_01334_),
    .B2(_04146_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09276_ (.A1(_01224_),
    .A2(_01232_),
    .A3(_01331_),
    .A4(_01333_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09277_ (.A1(_04181_),
    .A2(_04210_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(_01255_),
    .A2(_01339_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09279_ (.A1(_01247_),
    .A2(_04129_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09280_ (.A1(_04198_),
    .A2(_04212_),
    .A3(_04213_),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09281_ (.A1(_01226_),
    .A2(_01234_),
    .A3(net77),
    .A4(net76),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09282_ (.A1(_04209_),
    .A2(_04211_),
    .A3(_04214_),
    .B1(_04215_),
    .B2(_04182_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09283_ (.A1(_01255_),
    .A2(_04129_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09284_ (.A1(_01263_),
    .A2(_04131_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09285_ (.A1(_04171_),
    .A2(_04217_),
    .A3(_04218_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09286_ (.A1(_04182_),
    .A2(_04185_),
    .A3(_04219_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09287_ (.A1(_04216_),
    .A2(_04220_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09288_ (.A1(_04216_),
    .A2(_04220_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09289_ (.A1(_04208_),
    .A2(_04221_),
    .B(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09290_ (.A1(_04188_),
    .A2(_04189_),
    .A3(_04178_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09291_ (.A1(_04223_),
    .A2(_04224_),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09292_ (.A1(_04223_),
    .A2(_04224_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09293_ (.A1(_04206_),
    .A2(_04225_),
    .B(_04226_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09294_ (.A1(_04177_),
    .A2(_04194_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09295_ (.A1(_01227_),
    .A2(net74),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(_01243_),
    .A2(_01352_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09297_ (.A1(_01235_),
    .A2(_01348_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09298_ (.A1(_04230_),
    .A2(_04231_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09299_ (.A1(_04230_),
    .A2(_04231_),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09300_ (.A1(_04229_),
    .A2(_04232_),
    .B(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09301_ (.A1(_01242_),
    .A2(_01250_),
    .A3(_01347_),
    .A4(_01351_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09302_ (.A1(_01242_),
    .A2(_01347_),
    .B1(_01352_),
    .B2(_01250_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09303_ (.A1(_04235_),
    .A2(_04236_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09304_ (.A1(_01226_),
    .A2(_01234_),
    .A3(_04172_),
    .A4(_04169_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09305_ (.A1(_01226_),
    .A2(net75),
    .B1(net74),
    .B2(_01235_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09306_ (.A1(_04238_),
    .A2(_04239_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09307_ (.A1(_04237_),
    .A2(_04240_),
    .Z(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09308_ (.A1(_04234_),
    .A2(_04241_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09309_ (.A1(_04230_),
    .A2(_04231_),
    .A3(_04229_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09310_ (.A1(_01227_),
    .A2(_01235_),
    .A3(_01348_),
    .A4(_01353_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09311_ (.A1(_04243_),
    .A2(_04244_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09312_ (.A1(_04234_),
    .A2(_04241_),
    .Z(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09313_ (.A1(_04245_),
    .A2(_04246_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09314_ (.A1(_04242_),
    .A2(_04247_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(_01225_),
    .A2(_01335_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09316_ (.A1(_01242_),
    .A2(_01341_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09317_ (.A1(_01234_),
    .A2(_01338_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09318_ (.A1(_04249_),
    .A2(_04250_),
    .A3(_04251_),
    .Z(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09319_ (.A1(_01250_),
    .A2(_01346_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09320_ (.A1(_01258_),
    .A2(_01351_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09321_ (.A1(_04253_),
    .A2(_04238_),
    .A3(_04254_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09322_ (.A1(_04252_),
    .A2(_04255_),
    .Z(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09323_ (.A1(_04252_),
    .A2(_04255_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09324_ (.A1(_04256_),
    .A2(_04257_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09325_ (.A1(_04237_),
    .A2(_04240_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09326_ (.A1(_04235_),
    .A2(_04259_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09327_ (.A1(_04258_),
    .A2(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09328_ (.A1(_04258_),
    .A2(_04260_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09329_ (.A1(_04248_),
    .A2(_04261_),
    .B(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09330_ (.A1(_04253_),
    .A2(_04238_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09331_ (.A1(_04264_),
    .A2(_04254_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09332_ (.A1(_04253_),
    .A2(_04238_),
    .B(_04265_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09333_ (.A1(_01265_),
    .A2(_01350_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09334_ (.A1(_01232_),
    .A2(_04146_),
    .A3(_01337_),
    .A4(_04131_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09335_ (.A1(_01256_),
    .A2(_01346_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09336_ (.A1(_04268_),
    .A2(_04269_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09337_ (.A1(_04267_),
    .A2(_04270_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09338_ (.A1(_01241_),
    .A2(_01337_),
    .B1(_04131_),
    .B2(_01248_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09339_ (.A1(_01240_),
    .A2(_01247_),
    .A3(_01336_),
    .A4(_01340_),
    .Z(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09340_ (.I(_04273_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09341_ (.A1(_04272_),
    .A2(_04274_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09342_ (.A1(_01225_),
    .A2(_01332_),
    .B1(_01335_),
    .B2(_01233_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09343_ (.A1(_04210_),
    .A2(_04276_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09344_ (.A1(_01233_),
    .A2(_04172_),
    .B1(_04169_),
    .B2(_01241_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09345_ (.A1(_04249_),
    .A2(_04278_),
    .A3(_04268_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09346_ (.A1(_04275_),
    .A2(_04277_),
    .A3(_04279_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09347_ (.A1(_04271_),
    .A2(_04280_),
    .A3(_04256_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09348_ (.A1(_04266_),
    .A2(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09349_ (.A1(_04271_),
    .A2(_04280_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09350_ (.A1(_04256_),
    .A2(_04283_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09351_ (.A1(_04266_),
    .A2(_04281_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09352_ (.A1(_04284_),
    .A2(_04285_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09353_ (.A1(_04250_),
    .A2(_04251_),
    .A3(_04269_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09354_ (.A1(_04267_),
    .A2(_04270_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09355_ (.A1(_04287_),
    .A2(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09356_ (.A1(_01264_),
    .A2(_01345_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09357_ (.A1(_04273_),
    .A2(_04290_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09358_ (.A1(_01270_),
    .A2(_01351_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09359_ (.A1(_04291_),
    .A2(_04292_),
    .Z(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09360_ (.A1(_04209_),
    .A2(_04211_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09361_ (.A1(_04210_),
    .A2(_04272_),
    .A3(_04274_),
    .A4(_04276_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09362_ (.A1(_04294_),
    .A2(_04214_),
    .A3(_04295_),
    .Z(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09363_ (.A1(_04272_),
    .A2(_04274_),
    .B1(_04276_),
    .B2(_04210_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09364_ (.A1(_04295_),
    .A2(_04297_),
    .A3(_04279_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09365_ (.A1(_04271_),
    .A2(_04280_),
    .B(_04298_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09366_ (.A1(_04293_),
    .A2(_04296_),
    .A3(_04299_),
    .Z(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09367_ (.A1(_04289_),
    .A2(_04300_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09368_ (.A1(_04286_),
    .A2(_04301_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09369_ (.A1(_04263_),
    .A2(_04282_),
    .A3(_04302_),
    .B1(_04301_),
    .B2(_04286_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09370_ (.A1(_04293_),
    .A2(_04296_),
    .Z(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09371_ (.A1(_04293_),
    .A2(_04296_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09372_ (.A1(_04304_),
    .A2(_04299_),
    .A3(_04305_),
    .B1(_04289_),
    .B2(_04300_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09373_ (.A1(_01266_),
    .A2(_01348_),
    .A3(_04274_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09374_ (.A1(_04291_),
    .A2(_04292_),
    .B(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09375_ (.I(_04293_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09376_ (.A1(_04209_),
    .A2(_04211_),
    .A3(_04214_),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09377_ (.A1(_04209_),
    .A2(_04211_),
    .B(_04214_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09378_ (.A1(_04275_),
    .A2(_04277_),
    .Z(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09379_ (.A1(_04310_),
    .A2(_04311_),
    .B(_04312_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09380_ (.A1(_04310_),
    .A2(_04312_),
    .A3(_04311_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09381_ (.A1(_04309_),
    .A2(_04313_),
    .B(_04314_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09382_ (.A1(_04208_),
    .A2(_04221_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09383_ (.A1(_04315_),
    .A2(_04316_),
    .Z(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09384_ (.A1(_04308_),
    .A2(_04317_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09385_ (.A1(_04306_),
    .A2(_04318_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09386_ (.A1(_04306_),
    .A2(_04318_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09387_ (.A1(_04303_),
    .A2(_04319_),
    .B(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09388_ (.A1(_04315_),
    .A2(_04316_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09389_ (.A1(_04308_),
    .A2(_04317_),
    .B(_04322_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09390_ (.A1(_04206_),
    .A2(_04225_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09391_ (.A1(_04323_),
    .A2(_04324_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09392_ (.A1(_04323_),
    .A2(_04324_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09393_ (.A1(_04325_),
    .A2(_04326_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09394_ (.A1(_04321_),
    .A2(_04327_),
    .B(_04325_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09395_ (.A1(_04227_),
    .A2(_04228_),
    .Z(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09396_ (.A1(_04328_),
    .A2(_04329_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09397_ (.A1(_04227_),
    .A2(_04228_),
    .B(_04330_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09398_ (.A1(_04168_),
    .A2(_04196_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09399_ (.I(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09400_ (.A1(_04331_),
    .A2(_04333_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09401_ (.A1(_04197_),
    .A2(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09402_ (.A1(_04144_),
    .A2(_04165_),
    .Z(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09403_ (.A1(_04335_),
    .A2(_04336_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09404_ (.A1(_04166_),
    .A2(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09405_ (.A1(_04107_),
    .A2(_04093_),
    .A3(_04096_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09406_ (.A1(_04108_),
    .A2(_04339_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09407_ (.A1(_04119_),
    .A2(_04143_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09408_ (.A1(_04340_),
    .A2(_04341_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09409_ (.A1(_04340_),
    .A2(_04341_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09410_ (.A1(_04338_),
    .A2(_04342_),
    .B(_04343_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09411_ (.A1(_04108_),
    .A2(_04115_),
    .B1(_04118_),
    .B2(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09412_ (.I(_04112_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09413_ (.A1(_04346_),
    .A2(_04114_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09414_ (.A1(_04116_),
    .A2(_04115_),
    .B(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09415_ (.A1(_01975_),
    .A2(_04098_),
    .B1(_04109_),
    .B2(_04111_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09416_ (.A1(_01276_),
    .A2(_02081_),
    .A3(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09417_ (.A1(_04348_),
    .A2(_04350_),
    .Z(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09418_ (.A1(_01281_),
    .A2(net79),
    .A3(_04348_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09419_ (.A1(_04345_),
    .A2(_04351_),
    .B(_04352_),
    .C(_04349_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09420_ (.A1(_04059_),
    .A2(_04353_),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09421_ (.A1(_04345_),
    .A2(_04351_),
    .Z(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09422_ (.A1(_04344_),
    .A2(_04118_),
    .Z(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09423_ (.A1(_04338_),
    .A2(_04342_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09424_ (.A1(_04335_),
    .A2(_04336_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09425_ (.A1(_04331_),
    .A2(_04332_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09426_ (.A1(_04328_),
    .A2(_04329_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09427_ (.A1(_04321_),
    .A2(_04327_),
    .Z(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09428_ (.A1(_04306_),
    .A2(_04318_),
    .A3(_04303_),
    .Z(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09429_ (.A1(_04263_),
    .A2(_04282_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09430_ (.A1(_04363_),
    .A2(_04302_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09431_ (.A1(_04263_),
    .A2(_04282_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09432_ (.A1(_04363_),
    .A2(_04365_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09433_ (.A1(_04258_),
    .A2(_04260_),
    .A3(_04248_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09434_ (.A1(_04245_),
    .A2(_04246_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09435_ (.A1(_04243_),
    .A2(_04244_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09436_ (.A1(_01228_),
    .A2(net104),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09437_ (.A1(_01228_),
    .A2(net105),
    .B1(_01353_),
    .B2(_01236_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09438_ (.A1(_04368_),
    .A2(_04369_),
    .A3(_04370_),
    .A4(_04371_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09439_ (.A1(_04364_),
    .A2(_04366_),
    .A3(_04367_),
    .A4(_04372_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09440_ (.A1(_04360_),
    .A2(_04361_),
    .A3(_04362_),
    .A4(_04373_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09441_ (.A1(_04357_),
    .A2(_04358_),
    .A3(_04359_),
    .A4(_04374_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _09442_ (.A1(_04355_),
    .A2(_04356_),
    .A3(_04375_),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09443_ (.A1(_03819_),
    .A2(_03846_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09444_ (.A1(_03826_),
    .A2(_04058_),
    .B1(_04354_),
    .B2(_04376_),
    .C(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09445_ (.A1(_04005_),
    .A2(_04378_),
    .B(_03843_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09446_ (.A1(_01319_),
    .A2(_04004_),
    .B(_04379_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09447_ (.A1(_01084_),
    .A2(_03172_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09448_ (.A1(_03874_),
    .A2(_04009_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09449_ (.A1(_03875_),
    .A2(_04380_),
    .B(_04381_),
    .C(_04382_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _09450_ (.A1(_02228_),
    .A2(_01434_),
    .B1(_01457_),
    .B2(_02300_),
    .C1(_02929_),
    .C2(_01505_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09451_ (.A1(_02435_),
    .A2(_01492_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09452_ (.A1(_03274_),
    .A2(_03850_),
    .B1(_02420_),
    .B2(_02890_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09453_ (.A1(_02088_),
    .A2(_01101_),
    .B1(_01470_),
    .B2(_03060_),
    .C(_04386_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09454_ (.A1(_04381_),
    .A2(_04384_),
    .A3(_04385_),
    .A4(_04387_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09455_ (.A1(_03827_),
    .A2(_04388_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09456_ (.A1(_03993_),
    .A2(_04003_),
    .B1(_04383_),
    .B2(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09457_ (.I(_03821_),
    .Z(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09458_ (.A1(_04391_),
    .A2(_04380_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09459_ (.A1(_02930_),
    .A2(_03968_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(_02508_),
    .A2(_01319_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09461_ (.A1(_03883_),
    .A2(_04393_),
    .A3(_04394_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09462_ (.A1(_03895_),
    .A2(_04392_),
    .A3(_04395_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09463_ (.A1(_03896_),
    .A2(_04390_),
    .B(_04396_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09464_ (.A1(_03868_),
    .A2(_04397_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09465_ (.A1(_01289_),
    .A2(_02131_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09466_ (.I(_03882_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09467_ (.A1(_02622_),
    .A2(_04400_),
    .B(_03886_),
    .C(_02089_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09468_ (.A1(net67),
    .A2(_04391_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09469_ (.A1(_02930_),
    .A2(_01123_),
    .A3(_04402_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09470_ (.A1(\as2650.debug_psu[4] ),
    .A2(_04391_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09471_ (.A1(_02392_),
    .A2(_02189_),
    .A3(_04404_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09472_ (.I(_02597_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09473_ (.A1(_01579_),
    .A2(_03971_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09474_ (.A1(_04406_),
    .A2(_04400_),
    .B(_04407_),
    .C(_03061_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09475_ (.A1(_04401_),
    .A2(_04403_),
    .A3(_04405_),
    .A4(_04408_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09476_ (.A1(\as2650.debug_psu[7] ),
    .A2(_02186_),
    .B(_04025_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09477_ (.A1(_01569_),
    .A2(_04400_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09478_ (.A1(_01608_),
    .A2(_03897_),
    .B(_02834_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09479_ (.A1(_01573_),
    .A2(_03882_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09480_ (.A1(_02557_),
    .A2(_03971_),
    .B(_04413_),
    .C(_02301_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09481_ (.A1(_01629_),
    .A2(_03878_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09482_ (.A1(_01325_),
    .A2(_03878_),
    .B(_04415_),
    .C(_02435_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09483_ (.A1(_04414_),
    .A2(_04416_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09484_ (.A1(_02514_),
    .A2(_04410_),
    .B1(_04411_),
    .B2(_04412_),
    .C(_04417_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09485_ (.A1(_04409_),
    .A2(_04418_),
    .B(_03868_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09486_ (.A1(_03029_),
    .A2(_01289_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09487_ (.A1(_02180_),
    .A2(_02182_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09488_ (.A1(_04380_),
    .A2(_04399_),
    .B1(_04420_),
    .B2(_04421_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09489_ (.A1(_04398_),
    .A2(_04399_),
    .A3(_04419_),
    .B(_04422_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(_03993_),
    .A2(_04003_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09491_ (.A1(_04424_),
    .A2(_04382_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09492_ (.I(_02091_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09493_ (.A1(_04420_),
    .A2(_04425_),
    .B(_04426_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09494_ (.A1(_02947_),
    .A2(_02436_),
    .A3(_02392_),
    .A4(_03061_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09495_ (.A1(_03265_),
    .A2(_02835_),
    .A3(_03255_),
    .A4(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09496_ (.A1(_03274_),
    .A2(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09497_ (.I(_02939_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09498_ (.A1(_04423_),
    .A2(_04427_),
    .B1(_04430_),
    .B2(_04426_),
    .C(_04431_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09499_ (.A1(_04420_),
    .A2(_04421_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09500_ (.I(_04399_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09501_ (.A1(_01151_),
    .A2(_03843_),
    .A3(_03817_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _09502_ (.I(_02534_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09503_ (.A1(_03822_),
    .A2(_03820_),
    .A3(_03836_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09504_ (.A1(_04019_),
    .A2(_04410_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09505_ (.A1(_01326_),
    .A2(_04019_),
    .B(_04437_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09506_ (.A1(_03903_),
    .A2(_04438_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09507_ (.A1(_01280_),
    .A2(_03856_),
    .B1(_04436_),
    .B2(_01326_),
    .C(_04439_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09508_ (.A1(_03956_),
    .A2(_04440_),
    .B(_04016_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09509_ (.A1(_02543_),
    .A2(_04441_),
    .B(_04014_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09510_ (.A1(_04010_),
    .A2(_04442_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09511_ (.A1(_01281_),
    .A2(_04010_),
    .B(_03848_),
    .C(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09512_ (.A1(_04435_),
    .A2(_03848_),
    .B(_04444_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09513_ (.A1(_03829_),
    .A2(_04052_),
    .B(_03826_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09514_ (.A1(_03829_),
    .A2(_04445_),
    .B(_04446_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09515_ (.I(_03627_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09516_ (.A1(_04377_),
    .A2(_04354_),
    .A3(_04447_),
    .B1(_03847_),
    .B2(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09517_ (.A1(_01326_),
    .A2(_04434_),
    .B1(_04449_),
    .B2(_03844_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09518_ (.I(_04003_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09519_ (.A1(_03993_),
    .A2(_04451_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09520_ (.A1(_03874_),
    .A2(_02535_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09521_ (.A1(_03875_),
    .A2(_04450_),
    .B(_04453_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09522_ (.A1(_02180_),
    .A2(_04381_),
    .A3(_04454_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09523_ (.A1(_04452_),
    .A2(_04455_),
    .B(_03896_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09524_ (.A1(_02513_),
    .A2(_04024_),
    .B(_02188_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09525_ (.A1(_03888_),
    .A2(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09526_ (.A1(_02513_),
    .A2(_04025_),
    .B(_03881_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09527_ (.A1(_03897_),
    .A2(_04450_),
    .B1(_04458_),
    .B2(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09528_ (.A1(_04456_),
    .A2(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09529_ (.A1(_04433_),
    .A2(_04450_),
    .B1(_04461_),
    .B2(_03871_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09530_ (.A1(_02182_),
    .A2(_04435_),
    .B(_04452_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09531_ (.A1(_04432_),
    .A2(_04462_),
    .B1(_04463_),
    .B2(_04420_),
    .C(_04426_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09532_ (.A1(_03274_),
    .A2(_04426_),
    .B(_04464_),
    .C(_03893_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09533_ (.A1(_01849_),
    .A2(_03090_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09534_ (.I(_04465_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09535_ (.A1(_02187_),
    .A2(_01175_),
    .A3(_03898_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09536_ (.A1(_03895_),
    .A2(_04467_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09537_ (.A1(_01540_),
    .A2(_04468_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09538_ (.I(_04469_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09539_ (.I(_03888_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09540_ (.A1(_03255_),
    .A2(_01601_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09541_ (.A1(_03255_),
    .A2(_04471_),
    .B(_04472_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09542_ (.I(_03170_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09543_ (.I(_04474_),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09544_ (.I(_01857_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09545_ (.I(_03832_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09546_ (.A1(_03429_),
    .A2(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09547_ (.I(_04436_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09548_ (.A1(_01600_),
    .A2(_04436_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09549_ (.A1(_01854_),
    .A2(_04479_),
    .B(_04480_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09550_ (.A1(_04476_),
    .A2(_04478_),
    .A3(_04481_),
    .Z(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09551_ (.A1(_03257_),
    .A2(_04482_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09552_ (.A1(_01175_),
    .A2(_03179_),
    .A3(_01849_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09553_ (.A1(_01190_),
    .A2(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09554_ (.A1(_04468_),
    .A2(_04485_),
    .B(_03186_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09555_ (.A1(_02622_),
    .A2(_04475_),
    .B(_04483_),
    .C(_04486_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09556_ (.A1(_04470_),
    .A2(_04473_),
    .B(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09557_ (.A1(_01532_),
    .A2(_01190_),
    .A3(_04484_),
    .B(_04465_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09558_ (.A1(_04466_),
    .A2(_04488_),
    .B1(_04489_),
    .B2(_01601_),
    .C(_04431_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09559_ (.A1(_02625_),
    .A2(_02715_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09560_ (.I(_04469_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09561_ (.A1(_02228_),
    .A2(_02624_),
    .B(_03914_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09562_ (.I(_04476_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09563_ (.A1(_02594_),
    .A2(_02676_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09564_ (.I(_03173_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09565_ (.I(_04436_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09566_ (.A1(_01608_),
    .A2(_04479_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09567_ (.A1(_01898_),
    .A2(_04496_),
    .B(_04497_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09568_ (.A1(_01134_),
    .A2(_01126_),
    .A3(_04495_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09569_ (.A1(_04495_),
    .A2(_04498_),
    .B1(_04499_),
    .B2(_01608_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09570_ (.A1(_04494_),
    .A2(_04478_),
    .B1(_04500_),
    .B2(_04477_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09571_ (.A1(_04493_),
    .A2(_04490_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09572_ (.A1(_04493_),
    .A2(_04501_),
    .B(_04502_),
    .C(_04474_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09573_ (.A1(_02624_),
    .A2(_04475_),
    .B(_04486_),
    .C(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09574_ (.A1(_04491_),
    .A2(_04492_),
    .B(_04504_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09575_ (.A1(_04490_),
    .A2(_04489_),
    .B1(_04505_),
    .B2(_04466_),
    .C(_04431_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09576_ (.A1(_02596_),
    .A2(_02714_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09577_ (.A1(_00518_),
    .A2(_01615_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09578_ (.A1(_03265_),
    .A2(_04471_),
    .B(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09579_ (.A1(_02596_),
    .A2(_04479_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09580_ (.A1(_01914_),
    .A2(_04496_),
    .B(_04509_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09581_ (.A1(_01614_),
    .A2(_04499_),
    .B1(_04510_),
    .B2(_04495_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09582_ (.A1(_03156_),
    .A2(_04478_),
    .B1(_04511_),
    .B2(_04477_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09583_ (.A1(_04476_),
    .A2(_04506_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09584_ (.A1(_04493_),
    .A2(_04512_),
    .B(_04513_),
    .C(_04474_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09585_ (.A1(_02557_),
    .A2(_04475_),
    .B(_04486_),
    .C(_04514_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09586_ (.A1(_04491_),
    .A2(_04508_),
    .B(_04515_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09587_ (.A1(_04489_),
    .A2(_04506_),
    .B1(_04516_),
    .B2(_04466_),
    .C(_04431_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09588_ (.A1(_02556_),
    .A2(_02714_),
    .B(_02597_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09589_ (.A1(_02714_),
    .A2(_02677_),
    .B(_04517_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09590_ (.A1(_03062_),
    .A2(_04406_),
    .B(_03944_),
    .C(_04467_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09591_ (.A1(_01618_),
    .A2(_04479_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09592_ (.A1(_01928_),
    .A2(_04496_),
    .B(_04520_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09593_ (.A1(_02558_),
    .A2(_04499_),
    .B1(_04521_),
    .B2(_04495_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09594_ (.A1(_03139_),
    .A2(_04478_),
    .B1(_04522_),
    .B2(_04477_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09595_ (.A1(_04476_),
    .A2(_04518_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09596_ (.A1(_04493_),
    .A2(_04523_),
    .B(_04524_),
    .C(_04474_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09597_ (.A1(_04406_),
    .A2(_03260_),
    .B(_04486_),
    .C(_04525_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09598_ (.A1(_03750_),
    .A2(_04519_),
    .B(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09599_ (.A1(_04489_),
    .A2(_04518_),
    .B1(_04527_),
    .B2(_04466_),
    .C(_02987_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09600_ (.I(_03906_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09601_ (.I(_04496_),
    .Z(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09602_ (.A1(_04528_),
    .A2(_04529_),
    .B(_03040_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09603_ (.A1(_03793_),
    .A2(_04528_),
    .B1(_04529_),
    .B2(net100),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09604_ (.A1(_03258_),
    .A2(_04531_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09605_ (.A1(_01623_),
    .A2(_04530_),
    .B(_04532_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09606_ (.A1(_02890_),
    .A2(_01623_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09607_ (.A1(_03187_),
    .A2(_03951_),
    .A3(_04467_),
    .A4(_04534_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09608_ (.A1(_01184_),
    .A2(_04535_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09609_ (.A1(_04470_),
    .A2(_04533_),
    .B(_04536_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09610_ (.A1(_04400_),
    .A2(_03903_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09611_ (.A1(_01208_),
    .A2(_03176_),
    .B1(_04537_),
    .B2(_01962_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09612_ (.A1(_01630_),
    .A2(_04537_),
    .B1(_04538_),
    .B2(_03040_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09613_ (.A1(_03168_),
    .A2(_04528_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09614_ (.A1(_01630_),
    .A2(_03260_),
    .B(_04469_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09615_ (.A1(_04528_),
    .A2(_04539_),
    .B1(_04540_),
    .B2(_03258_),
    .C(_04541_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09616_ (.A1(_02436_),
    .A2(_01630_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09617_ (.A1(_02437_),
    .A2(_04471_),
    .B(_04491_),
    .C(_04543_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09618_ (.A1(_02987_),
    .A2(_04542_),
    .A3(_04544_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09619_ (.I(_04545_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09620_ (.A1(_03207_),
    .A2(_03906_),
    .B1(_04529_),
    .B2(net102),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09621_ (.A1(_04475_),
    .A2(_04546_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09622_ (.A1(_01633_),
    .A2(_04530_),
    .B(_04547_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09623_ (.I(_04491_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09624_ (.A1(_02508_),
    .A2(_01633_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09625_ (.A1(_04393_),
    .A2(_04549_),
    .A3(_04550_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09626_ (.A1(_04470_),
    .A2(_04548_),
    .B(_04551_),
    .C(_03893_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09627_ (.A1(_03252_),
    .A2(_03907_),
    .B1(_04529_),
    .B2(net103),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09628_ (.A1(_03910_),
    .A2(_04552_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09629_ (.A1(net5),
    .A2(_04530_),
    .B(_04553_),
    .C(_04470_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09630_ (.A1(_03071_),
    .A2(_04471_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09631_ (.A1(_03071_),
    .A2(_01636_),
    .B(_04549_),
    .C(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09632_ (.A1(_04554_),
    .A2(_04556_),
    .B(_01529_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09633_ (.A1(_01399_),
    .A2(_01412_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09634_ (.A1(_02179_),
    .A2(_02187_),
    .B(_03921_),
    .C(_00505_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09635_ (.A1(_02179_),
    .A2(_03887_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09636_ (.A1(_02213_),
    .A2(_04557_),
    .A3(_04558_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09637_ (.I(_04559_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09638_ (.I(_04560_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09639_ (.I(_02169_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09640_ (.I(_01437_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09641_ (.A1(_01947_),
    .A2(_02219_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09642_ (.I(_04564_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09643_ (.A1(_04563_),
    .A2(_04565_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09644_ (.A1(_01856_),
    .A2(_02197_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09645_ (.A1(_03816_),
    .A2(_04567_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09646_ (.A1(_01134_),
    .A2(_01393_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09647_ (.A1(_04569_),
    .A2(_04567_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09648_ (.I(_01862_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09649_ (.A1(_03833_),
    .A2(_03825_),
    .B(_04571_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09650_ (.A1(_01863_),
    .A2(_03838_),
    .A3(_03813_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09651_ (.A1(_01394_),
    .A2(_04571_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09652_ (.A1(_04573_),
    .A2(_04574_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09653_ (.A1(_04568_),
    .A2(_04570_),
    .A3(_04572_),
    .A4(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09654_ (.I(_04576_),
    .Z(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09655_ (.A1(_04566_),
    .A2(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09656_ (.I(_04578_),
    .Z(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09657_ (.A1(_01361_),
    .A2(\as2650.regs[4][0] ),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09658_ (.A1(_00650_),
    .A2(_02207_),
    .Z(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09659_ (.A1(_04563_),
    .A2(_04581_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09660_ (.A1(_01181_),
    .A2(_04582_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09661_ (.I(_04583_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09662_ (.I(_04584_),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09663_ (.I(_04568_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09664_ (.I(_04586_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09665_ (.A1(_04569_),
    .A2(_04567_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09666_ (.I(_04588_),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09667_ (.I(_04589_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09668_ (.I(_04573_),
    .Z(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09669_ (.I(_04591_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09670_ (.A1(_01394_),
    .A2(_01863_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09671_ (.I(_04593_),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09672_ (.A1(_01856_),
    .A2(_02198_),
    .A3(_03832_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09673_ (.I(_04595_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09674_ (.A1(_03331_),
    .A2(_04595_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09675_ (.A1(_02002_),
    .A2(_04596_),
    .B(_04597_),
    .C(_04593_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09676_ (.A1(_04571_),
    .A2(_04059_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09677_ (.I(_04599_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09678_ (.A1(\as2650.chirpchar[0] ),
    .A2(_04594_),
    .B(_04598_),
    .C(_04600_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09679_ (.A1(_02198_),
    .A2(_03826_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09680_ (.I(_04602_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09681_ (.A1(net73),
    .A2(net104),
    .A3(_04603_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09682_ (.I(_04591_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09683_ (.A1(_04601_),
    .A2(_04604_),
    .B(_04605_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09684_ (.A1(_02126_),
    .A2(_04592_),
    .B(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09685_ (.A1(_01556_),
    .A2(_04589_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09686_ (.I(_04586_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09687_ (.A1(_04590_),
    .A2(_04607_),
    .B(_04608_),
    .C(_04609_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09688_ (.A1(_01601_),
    .A2(_04587_),
    .B(_04610_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09689_ (.A1(_03947_),
    .A2(_04577_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09690_ (.I(_04612_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09691_ (.A1(_04580_),
    .A2(_04585_),
    .B1(_04611_),
    .B2(_04613_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09692_ (.A1(_04562_),
    .A2(_04579_),
    .B(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09693_ (.I(_04560_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09694_ (.A1(_01948_),
    .A2(_04559_),
    .A3(_04583_),
    .A4(_04577_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09695_ (.I(_04617_),
    .Z(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09696_ (.A1(_02211_),
    .A2(_04616_),
    .B1(_04618_),
    .B2(\as2650.regs[0][0] ),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09697_ (.A1(_04561_),
    .A2(_04615_),
    .B(_04619_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09698_ (.A1(_02835_),
    .A2(_02384_),
    .B1(_02289_),
    .B2(_02292_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09699_ (.A1(_01361_),
    .A2(\as2650.regs[4][1] ),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09700_ (.I(_04586_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09701_ (.A1(_04571_),
    .A2(_03838_),
    .A3(_03815_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09702_ (.I(_04371_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09703_ (.A1(_04244_),
    .A2(_04624_),
    .B(_04600_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09704_ (.A1(_03845_),
    .A2(_04567_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09705_ (.I(_04626_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09706_ (.A1(_03381_),
    .A2(_04627_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09707_ (.A1(_02016_),
    .A2(_04627_),
    .B(_04628_),
    .C(_04574_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09708_ (.I(_04602_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09709_ (.A1(\as2650.chirpchar[1] ),
    .A2(_04574_),
    .B(_04629_),
    .C(_04630_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09710_ (.A1(_04625_),
    .A2(_04631_),
    .B(_04623_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09711_ (.A1(_02266_),
    .A2(_04623_),
    .B(_04632_),
    .C(_04570_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09712_ (.I(_04586_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09713_ (.A1(_03901_),
    .A2(_04570_),
    .B(_04633_),
    .C(_04634_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09714_ (.A1(_01609_),
    .A2(_04622_),
    .B(_04635_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09715_ (.A1(_04621_),
    .A2(_04585_),
    .B1(_04613_),
    .B2(_04636_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09716_ (.A1(_04620_),
    .A2(_04579_),
    .B(_04637_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09717_ (.I(_02266_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09718_ (.I(_04559_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09719_ (.A1(_04639_),
    .A2(_04640_),
    .B1(_04618_),
    .B2(\as2650.regs[0][1] ),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09720_ (.A1(_04561_),
    .A2(_04638_),
    .B(_04641_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09721_ (.A1(_03265_),
    .A2(_02384_),
    .B1(_02337_),
    .B2(_02338_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09722_ (.A1(_01361_),
    .A2(\as2650.regs[4][2] ),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09723_ (.I(_04589_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09724_ (.I(_04591_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09725_ (.I(_04630_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09726_ (.I(_04627_),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09727_ (.I(_04626_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09728_ (.A1(_02031_),
    .A2(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09729_ (.A1(_03427_),
    .A2(_04647_),
    .B(_04649_),
    .C(_04594_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09730_ (.I(_04574_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09731_ (.A1(\as2650.chirpchar[2] ),
    .A2(_04651_),
    .B(_04603_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09732_ (.A1(_04369_),
    .A2(_04646_),
    .B1(_04650_),
    .B2(_04652_),
    .C(_04605_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09733_ (.A1(_02326_),
    .A2(_04645_),
    .B(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09734_ (.I(_04588_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09735_ (.A1(_01574_),
    .A2(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09736_ (.A1(_04644_),
    .A2(_04654_),
    .B(_04656_),
    .C(_04634_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09737_ (.A1(_01615_),
    .A2(_04622_),
    .B(_04657_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09738_ (.A1(_04643_),
    .A2(_04585_),
    .B1(_04613_),
    .B2(_04658_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09739_ (.A1(_04642_),
    .A2(_04579_),
    .B(_04659_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09740_ (.I(_02326_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09741_ (.A1(_04661_),
    .A2(_04640_),
    .B1(_04618_),
    .B2(\as2650.regs[0][2] ),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09742_ (.A1(_04561_),
    .A2(_04660_),
    .B(_04662_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09743_ (.A1(_02385_),
    .A2(_02382_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09744_ (.I(_01360_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09745_ (.A1(_04664_),
    .A2(\as2650.regs[4][3] ),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09746_ (.I(_04612_),
    .Z(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09747_ (.I(_04627_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09748_ (.A1(_02044_),
    .A2(_04648_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09749_ (.A1(_03469_),
    .A2(_04667_),
    .B(_04668_),
    .C(_04594_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09750_ (.A1(\as2650.chirpchar[3] ),
    .A2(_04651_),
    .B(_04603_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09751_ (.A1(_04368_),
    .A2(_04646_),
    .B1(_04669_),
    .B2(_04670_),
    .C(_04605_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09752_ (.A1(_02369_),
    .A2(_04645_),
    .B(_04671_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09753_ (.A1(_01579_),
    .A2(_04655_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09754_ (.A1(_04644_),
    .A2(_04672_),
    .B(_04673_),
    .C(_04634_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09755_ (.A1(_01619_),
    .A2(_04622_),
    .B(_04674_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09756_ (.A1(_04665_),
    .A2(_04585_),
    .B1(_04666_),
    .B2(_04675_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09757_ (.A1(_04663_),
    .A2(_04579_),
    .B(_04676_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09758_ (.I(_02369_),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09759_ (.A1(_04678_),
    .A2(_04640_),
    .B1(_04618_),
    .B2(\as2650.regs[0][3] ),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09760_ (.A1(_04561_),
    .A2(_04677_),
    .B(_04679_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09761_ (.I(_02430_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09762_ (.A1(_04664_),
    .A2(\as2650.regs[4][4] ),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09763_ (.A1(_03510_),
    .A2(_04595_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09764_ (.I(_04593_),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09765_ (.A1(_02054_),
    .A2(_04596_),
    .B(_04682_),
    .C(_04683_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09766_ (.A1(\as2650.chirpchar[4] ),
    .A2(_04594_),
    .B(_04684_),
    .C(_04600_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09767_ (.A1(_04367_),
    .A2(_04599_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09768_ (.A1(_04685_),
    .A2(_04686_),
    .B(_04592_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09769_ (.A1(_02419_),
    .A2(_04645_),
    .B(_04687_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09770_ (.A1(_01948_),
    .A2(_04655_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09771_ (.A1(_04644_),
    .A2(_04688_),
    .B(_04689_),
    .C(_04609_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09772_ (.A1(_01623_),
    .A2(_04587_),
    .B(_04690_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09773_ (.A1(_04681_),
    .A2(_04584_),
    .B1(_04666_),
    .B2(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09774_ (.A1(_04680_),
    .A2(_04578_),
    .B(_04692_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09775_ (.I(_02419_),
    .Z(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09776_ (.A1(_04694_),
    .A2(_04640_),
    .B1(_04617_),
    .B2(\as2650.regs[0][4] ),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09777_ (.A1(_04616_),
    .A2(_04693_),
    .B(_04695_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09778_ (.A1(_02915_),
    .A2(_02384_),
    .B1(_02468_),
    .B2(_02470_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09779_ (.A1(_04664_),
    .A2(\as2650.regs[4][5] ),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09780_ (.A1(_02067_),
    .A2(_04648_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09781_ (.A1(_03552_),
    .A2(_04667_),
    .B(_04698_),
    .C(_04683_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09782_ (.A1(\as2650.chirpchar[5] ),
    .A2(_04651_),
    .B(_04630_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09783_ (.A1(_04366_),
    .A2(_04646_),
    .B1(_04699_),
    .B2(_04700_),
    .C(_04605_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09784_ (.A1(_02458_),
    .A2(_04645_),
    .B(_04701_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09785_ (.A1(_01592_),
    .A2(_04655_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09786_ (.A1(_04590_),
    .A2(_04702_),
    .B(_04703_),
    .C(_04609_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09787_ (.A1(_01629_),
    .A2(_04587_),
    .B(_04704_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09788_ (.A1(_04697_),
    .A2(_04584_),
    .B1(_04666_),
    .B2(_04705_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09789_ (.A1(_04696_),
    .A2(_04578_),
    .B(_04706_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09790_ (.I(_02458_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09791_ (.A1(_04708_),
    .A2(_04560_),
    .B1(_04617_),
    .B2(\as2650.regs[0][5] ),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09792_ (.A1(_04616_),
    .A2(_04707_),
    .B(_04709_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09793_ (.A1(_02507_),
    .A2(_02509_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09794_ (.A1(_04664_),
    .A2(\as2650.regs[4][6] ),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09795_ (.A1(_02074_),
    .A2(_04648_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09796_ (.A1(_03593_),
    .A2(_04667_),
    .B(_04712_),
    .C(_04683_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09797_ (.A1(\as2650.chirpchar[6] ),
    .A2(_04651_),
    .B(_04630_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09798_ (.A1(_04364_),
    .A2(_04646_),
    .B1(_04713_),
    .B2(_04714_),
    .C(_04591_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09799_ (.A1(_02494_),
    .A2(_04592_),
    .B(_04715_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09800_ (.A1(_01320_),
    .A2(_04589_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09801_ (.A1(_04590_),
    .A2(_04716_),
    .B(_04717_),
    .C(_04609_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09802_ (.A1(_01633_),
    .A2(_04587_),
    .B(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09803_ (.A1(_04711_),
    .A2(_04584_),
    .B1(_04666_),
    .B2(_04719_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09804_ (.A1(_04710_),
    .A2(_04578_),
    .B(_04720_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09805_ (.I(_02494_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09806_ (.A1(_04722_),
    .A2(_04560_),
    .B1(_04617_),
    .B2(\as2650.regs[0][6] ),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09807_ (.A1(_04616_),
    .A2(_04721_),
    .B(_04723_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09808_ (.A1(_03948_),
    .A2(_04557_),
    .A3(_04558_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09809_ (.I(_04599_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09810_ (.A1(net79),
    .A2(_04596_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09811_ (.A1(_03627_),
    .A2(_04667_),
    .B(_04683_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09812_ (.A1(_04726_),
    .A2(_04727_),
    .B(_04600_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09813_ (.A1(_04362_),
    .A2(_04725_),
    .B(_04728_),
    .C(_04623_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09814_ (.A1(_02554_),
    .A2(_04592_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09815_ (.A1(_04729_),
    .A2(_04730_),
    .B(_04590_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09816_ (.A1(_01327_),
    .A2(_04644_),
    .B(_04731_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09817_ (.A1(_01636_),
    .A2(_04634_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09818_ (.A1(_04622_),
    .A2(_04732_),
    .B(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09819_ (.A1(_01302_),
    .A2(net103),
    .A3(_04566_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09820_ (.A1(_02552_),
    .A2(_04582_),
    .B(_04612_),
    .C(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09821_ (.A1(_04613_),
    .A2(_04734_),
    .B(_04736_),
    .C(_04724_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09822_ (.A1(_04435_),
    .A2(_04724_),
    .B(_04737_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09823_ (.A1(_02178_),
    .A2(_03883_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09824_ (.I(_01947_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09825_ (.A1(_04739_),
    .A2(_02178_),
    .A3(_03883_),
    .A4(_02185_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09826_ (.I(_04740_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09827_ (.A1(_04738_),
    .A2(_04581_),
    .A3(_04741_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09828_ (.I(_04742_),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09829_ (.I(_04740_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09830_ (.A1(_04738_),
    .A2(_04565_),
    .B(_04740_),
    .C(_02222_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09831_ (.I(_04745_),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09832_ (.A1(_02211_),
    .A2(_04744_),
    .B1(_04746_),
    .B2(\as2650.regs[2][0] ),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09833_ (.A1(_02170_),
    .A2(_04743_),
    .B(_04747_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09834_ (.A1(_04639_),
    .A2(_04744_),
    .B1(_04746_),
    .B2(\as2650.regs[2][1] ),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09835_ (.A1(_02294_),
    .A2(_04743_),
    .B(_04748_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09836_ (.A1(_04661_),
    .A2(_04744_),
    .B1(_04746_),
    .B2(\as2650.regs[2][2] ),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09837_ (.A1(_02340_),
    .A2(_04743_),
    .B(_04749_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09838_ (.A1(_04678_),
    .A2(_04744_),
    .B1(_04746_),
    .B2(\as2650.regs[2][3] ),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09839_ (.A1(_02386_),
    .A2(_04743_),
    .B(_04750_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09840_ (.I(_04742_),
    .Z(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09841_ (.I(_04740_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09842_ (.I(_04745_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09843_ (.A1(_04694_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\as2650.regs[2][4] ),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09844_ (.A1(_02431_),
    .A2(_04751_),
    .B(_04754_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09845_ (.A1(_04708_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\as2650.regs[2][5] ),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09846_ (.A1(_02472_),
    .A2(_04751_),
    .B(_04755_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09847_ (.A1(_04722_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\as2650.regs[2][6] ),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09848_ (.A1(_02510_),
    .A2(_04751_),
    .B(_04756_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09849_ (.I(_02554_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09850_ (.A1(_04757_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\as2650.regs[2][7] ),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09851_ (.A1(_02553_),
    .A2(_04751_),
    .B(_04758_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09852_ (.I(_01413_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09853_ (.A1(_02213_),
    .A2(_03831_),
    .A3(_02185_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09854_ (.I(_04759_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09855_ (.I(_04760_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09856_ (.I(_04572_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09857_ (.A1(_03947_),
    .A2(_04762_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09858_ (.I(_04763_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09859_ (.I(_04603_),
    .Z(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09860_ (.I(_04765_),
    .Z(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09861_ (.A1(_04361_),
    .A2(_04766_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09862_ (.I(_04647_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09863_ (.A1(_01854_),
    .A2(_04647_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09864_ (.A1(_03654_),
    .A2(_04768_),
    .B(_04769_),
    .C(_04725_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09865_ (.A1(_04767_),
    .A2(_04770_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09866_ (.I(_03835_),
    .Z(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09867_ (.A1(_04772_),
    .A2(_02221_),
    .A3(_04762_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09868_ (.I(_04773_),
    .Z(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09869_ (.A1(_04764_),
    .A2(_04771_),
    .B1(_04774_),
    .B2(_04562_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09870_ (.I(_04760_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09871_ (.A1(_00507_),
    .A2(_04759_),
    .A3(_04763_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09872_ (.A1(_04772_),
    .A2(_02221_),
    .B(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09873_ (.I(_04778_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09874_ (.A1(_02211_),
    .A2(_04776_),
    .B1(_04779_),
    .B2(\as2650.regs[5][0] ),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09875_ (.A1(_04761_),
    .A2(_04775_),
    .B(_04780_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09876_ (.I(_04765_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09877_ (.I(_04647_),
    .Z(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09878_ (.A1(_01898_),
    .A2(_04782_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09879_ (.A1(_03702_),
    .A2(_04768_),
    .B(_04783_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09880_ (.A1(_04360_),
    .A2(_04766_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09881_ (.A1(_04781_),
    .A2(_04784_),
    .B(_04785_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09882_ (.I(_04764_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09883_ (.A1(_04620_),
    .A2(_04774_),
    .B1(_04786_),
    .B2(_04787_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09884_ (.A1(_04639_),
    .A2(_04776_),
    .B1(_04779_),
    .B2(\as2650.regs[5][1] ),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09885_ (.A1(_04761_),
    .A2(_04788_),
    .B(_04789_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09886_ (.I(_04596_),
    .Z(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09887_ (.I(_04790_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09888_ (.A1(_01914_),
    .A2(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09889_ (.I(_04765_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09890_ (.A1(_03727_),
    .A2(_04791_),
    .B(_04792_),
    .C(_04793_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09891_ (.A1(_04359_),
    .A2(_04781_),
    .B(_04794_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09892_ (.A1(_04642_),
    .A2(_04774_),
    .B1(_04795_),
    .B2(_04787_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09893_ (.A1(_04661_),
    .A2(_04776_),
    .B1(_04779_),
    .B2(\as2650.regs[5][2] ),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09894_ (.A1(_04761_),
    .A2(_04796_),
    .B(_04797_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09895_ (.A1(_03766_),
    .A2(_04791_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09896_ (.A1(net99),
    .A2(_04782_),
    .B(_04798_),
    .C(_04793_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09897_ (.A1(_04358_),
    .A2(_04781_),
    .B(_04799_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09898_ (.A1(_04663_),
    .A2(_04774_),
    .B1(_04800_),
    .B2(_04787_),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09899_ (.A1(_04678_),
    .A2(_04776_),
    .B1(_04779_),
    .B2(\as2650.regs[5][3] ),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09900_ (.A1(_04761_),
    .A2(_04801_),
    .B(_04802_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09901_ (.I(_04760_),
    .Z(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09902_ (.I(_04773_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09903_ (.A1(_03793_),
    .A2(_04790_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09904_ (.A1(net100),
    .A2(_04782_),
    .B(_04805_),
    .C(_04793_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09905_ (.A1(_04357_),
    .A2(_04781_),
    .B(_04806_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09906_ (.A1(_04680_),
    .A2(_04804_),
    .B1(_04807_),
    .B2(_04787_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09907_ (.I(_04760_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09908_ (.I(_04778_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09909_ (.A1(_04694_),
    .A2(_04809_),
    .B1(_04810_),
    .B2(\as2650.regs[5][4] ),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09910_ (.A1(_04803_),
    .A2(_04808_),
    .B(_04811_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09911_ (.A1(_04356_),
    .A2(_04766_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09912_ (.A1(_01962_),
    .A2(_04782_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09913_ (.A1(_03168_),
    .A2(_04768_),
    .B(_04813_),
    .C(_04725_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09914_ (.A1(_04812_),
    .A2(_04814_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09915_ (.A1(_04696_),
    .A2(_04804_),
    .B1(_04815_),
    .B2(_04764_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09916_ (.A1(_04708_),
    .A2(_04809_),
    .B1(_04810_),
    .B2(\as2650.regs[5][5] ),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09917_ (.A1(_04803_),
    .A2(_04816_),
    .B(_04817_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09918_ (.A1(_03207_),
    .A2(_04768_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09919_ (.A1(net102),
    .A2(_04791_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09920_ (.A1(_04355_),
    .A2(_04793_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09921_ (.A1(_04766_),
    .A2(_04818_),
    .A3(_04819_),
    .B(_04820_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09922_ (.A1(_04710_),
    .A2(_04804_),
    .B1(_04821_),
    .B2(_04764_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09923_ (.A1(_04722_),
    .A2(_04809_),
    .B1(_04810_),
    .B2(\as2650.regs[5][6] ),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09924_ (.A1(_04803_),
    .A2(_04822_),
    .B(_04823_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09925_ (.A1(_03252_),
    .A2(_04790_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09926_ (.A1(_01987_),
    .A2(_04790_),
    .B(_04824_),
    .C(_04725_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09927_ (.A1(_04353_),
    .A2(_04765_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09928_ (.A1(_04825_),
    .A2(_04826_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09929_ (.I(_04804_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09930_ (.A1(_03948_),
    .A2(_04762_),
    .A3(_04827_),
    .B1(_04828_),
    .B2(_02552_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09931_ (.I(_04829_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09932_ (.A1(_04757_),
    .A2(_04809_),
    .B1(_04810_),
    .B2(\as2650.regs[5][7] ),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09933_ (.A1(_04803_),
    .A2(_04830_),
    .B(_04831_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09934_ (.A1(_01358_),
    .A2(_03831_),
    .A3(_02184_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09935_ (.I(_04832_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09936_ (.I(_04833_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09937_ (.I(_04834_),
    .Z(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09938_ (.A1(_01947_),
    .A2(_04572_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09939_ (.I(_04836_),
    .Z(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09940_ (.A1(_04772_),
    .A2(_04564_),
    .A3(_04762_),
    .Z(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09941_ (.I(_04838_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09942_ (.A1(_04771_),
    .A2(_04837_),
    .B1(_04839_),
    .B2(_04562_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09943_ (.I(_02126_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09944_ (.I(_04833_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09945_ (.A1(_00506_),
    .A2(_04832_),
    .A3(_04836_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09946_ (.A1(_04772_),
    .A2(_04565_),
    .B(_04843_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09947_ (.I(_04844_),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09948_ (.A1(_04841_),
    .A2(_04842_),
    .B1(_04845_),
    .B2(\as2650.regs[1][0] ),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09949_ (.A1(_04835_),
    .A2(_04840_),
    .B(_04846_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09950_ (.A1(_04786_),
    .A2(_04837_),
    .B1(_04839_),
    .B2(_04620_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09951_ (.I(_04833_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09952_ (.A1(_04639_),
    .A2(_04848_),
    .B1(_04845_),
    .B2(\as2650.regs[1][1] ),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09953_ (.A1(_04835_),
    .A2(_04847_),
    .B(_04849_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09954_ (.A1(_04795_),
    .A2(_04837_),
    .B1(_04839_),
    .B2(_04642_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09955_ (.A1(_04661_),
    .A2(_04848_),
    .B1(_04845_),
    .B2(\as2650.regs[1][2] ),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09956_ (.A1(_04835_),
    .A2(_04850_),
    .B(_04851_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09957_ (.A1(_04800_),
    .A2(_04837_),
    .B1(_04839_),
    .B2(_04663_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09958_ (.A1(_04678_),
    .A2(_04848_),
    .B1(_04845_),
    .B2(\as2650.regs[1][3] ),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09959_ (.A1(_04835_),
    .A2(_04852_),
    .B(_04853_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09960_ (.I(_04836_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09961_ (.I(_04838_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09962_ (.A1(_04807_),
    .A2(_04854_),
    .B1(_04855_),
    .B2(_04680_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09963_ (.I(_04844_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09964_ (.A1(_04694_),
    .A2(_04848_),
    .B1(_04857_),
    .B2(\as2650.regs[1][4] ),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09965_ (.A1(_04842_),
    .A2(_04856_),
    .B(_04858_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09966_ (.A1(_04815_),
    .A2(_04854_),
    .B1(_04855_),
    .B2(_04696_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09967_ (.A1(_04708_),
    .A2(_04834_),
    .B1(_04857_),
    .B2(\as2650.regs[1][5] ),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09968_ (.A1(_04842_),
    .A2(_04859_),
    .B(_04860_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09969_ (.A1(_04821_),
    .A2(_04854_),
    .B1(_04855_),
    .B2(_04710_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09970_ (.A1(_04722_),
    .A2(_04834_),
    .B1(_04857_),
    .B2(\as2650.regs[1][6] ),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09971_ (.A1(_04842_),
    .A2(_04861_),
    .B(_04862_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09972_ (.I(_04827_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09973_ (.A1(_04863_),
    .A2(_04854_),
    .B(_04833_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09974_ (.A1(_02514_),
    .A2(_02230_),
    .B(_02551_),
    .C(_04855_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09975_ (.A1(_04435_),
    .A2(_04834_),
    .B1(_04864_),
    .B2(_04865_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09976_ (.I0(_04866_),
    .I1(\as2650.regs[1][7] ),
    .S(_04857_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09977_ (.I(_04867_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09978_ (.A1(_04739_),
    .A2(_04557_),
    .A3(_04558_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09979_ (.I(_04868_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09980_ (.I(_04869_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09981_ (.A1(_03947_),
    .A2(_01202_),
    .A3(_02219_),
    .A4(_04577_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09982_ (.I(_04871_),
    .Z(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09983_ (.A1(_01359_),
    .A2(_04576_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09984_ (.I(_04873_),
    .Z(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09985_ (.A1(_04563_),
    .A2(_02220_),
    .B(_00506_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09986_ (.I(_04875_),
    .Z(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09987_ (.A1(_01221_),
    .A2(_04876_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09988_ (.A1(_04611_),
    .A2(_04874_),
    .B(_04877_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09989_ (.A1(_04562_),
    .A2(_04872_),
    .B(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09990_ (.I(_04869_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09991_ (.I(_04576_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09992_ (.A1(_04739_),
    .A2(_04557_),
    .A3(_04558_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09993_ (.I(_04875_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09994_ (.A1(_01360_),
    .A2(_04881_),
    .A3(_04882_),
    .A4(_04883_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09995_ (.I(_04884_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09996_ (.A1(_04841_),
    .A2(_04880_),
    .B1(_04885_),
    .B2(\as2650.regs[4][0] ),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09997_ (.A1(_04870_),
    .A2(_04879_),
    .B(_04886_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09998_ (.A1(_01229_),
    .A2(_04876_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09999_ (.A1(_04636_),
    .A2(_04874_),
    .B(_04887_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10000_ (.A1(_04620_),
    .A2(_04872_),
    .B(_04888_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10001_ (.I(_04868_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10002_ (.A1(_02296_),
    .A2(_04890_),
    .B1(_04885_),
    .B2(\as2650.regs[4][1] ),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10003_ (.A1(_04870_),
    .A2(_04889_),
    .B(_04891_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10004_ (.A1(_01237_),
    .A2(_04876_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10005_ (.A1(_04658_),
    .A2(_04874_),
    .B(_04892_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10006_ (.A1(_04642_),
    .A2(_04872_),
    .B(_04893_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10007_ (.A1(_02341_),
    .A2(_04890_),
    .B1(_04885_),
    .B2(\as2650.regs[4][2] ),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10008_ (.A1(_04870_),
    .A2(_04894_),
    .B(_04895_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10009_ (.A1(_01245_),
    .A2(_04876_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10010_ (.A1(_04675_),
    .A2(_04874_),
    .B(_04896_),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10011_ (.A1(_04663_),
    .A2(_04872_),
    .B(_04897_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10012_ (.A1(_02387_),
    .A2(_04890_),
    .B1(_04885_),
    .B2(\as2650.regs[4][3] ),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10013_ (.A1(_04870_),
    .A2(_04898_),
    .B(_04899_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10014_ (.I(_04873_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10015_ (.A1(_01252_),
    .A2(_04883_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10016_ (.A1(_04691_),
    .A2(_04900_),
    .B(_04901_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10017_ (.A1(_04680_),
    .A2(_04871_),
    .B(_04902_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10018_ (.A1(_02432_),
    .A2(_04890_),
    .B1(_04884_),
    .B2(\as2650.regs[4][4] ),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10019_ (.A1(_04880_),
    .A2(_04903_),
    .B(_04904_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10020_ (.A1(_01260_),
    .A2(_04883_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10021_ (.A1(_04705_),
    .A2(_04900_),
    .B(_04905_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10022_ (.A1(_04696_),
    .A2(_04871_),
    .B(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10023_ (.A1(_02473_),
    .A2(_04869_),
    .B1(_04884_),
    .B2(\as2650.regs[4][5] ),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10024_ (.A1(_04880_),
    .A2(_04907_),
    .B(_04908_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10025_ (.A1(_01267_),
    .A2(_04883_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10026_ (.A1(_04719_),
    .A2(_04900_),
    .B(_04909_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10027_ (.A1(_04710_),
    .A2(_04871_),
    .B(_04910_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10028_ (.A1(_02511_),
    .A2(_04869_),
    .B1(_04884_),
    .B2(\as2650.regs[4][6] ),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10029_ (.A1(_04880_),
    .A2(_04911_),
    .B(_04912_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10030_ (.A1(_04563_),
    .A2(_02208_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10031_ (.A1(_01182_),
    .A2(net103),
    .A3(_04913_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10032_ (.A1(_02552_),
    .A2(_04913_),
    .B(_04914_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10033_ (.I0(_04734_),
    .I1(_04915_),
    .S(_04900_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10034_ (.I0(_04757_),
    .I1(_04916_),
    .S(_04882_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10035_ (.I(_04917_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10036_ (.I(_02185_),
    .Z(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10037_ (.A1(_02176_),
    .A2(_04918_),
    .A3(_04581_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10038_ (.I(_04919_),
    .Z(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10039_ (.A1(_01948_),
    .A2(_02178_),
    .A3(_04391_),
    .A4(_04918_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10040_ (.I(_04921_),
    .Z(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10041_ (.A1(_02176_),
    .A2(_04565_),
    .B(_04921_),
    .C(_02222_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10042_ (.I(_04923_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10043_ (.A1(_04841_),
    .A2(_04922_),
    .B1(_04924_),
    .B2(\as2650.regs[3][0] ),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10044_ (.A1(_02170_),
    .A2(_04920_),
    .B(_04925_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10045_ (.A1(_02296_),
    .A2(_04922_),
    .B1(_04924_),
    .B2(\as2650.regs[3][1] ),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10046_ (.A1(_02294_),
    .A2(_04920_),
    .B(_04926_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10047_ (.A1(_02341_),
    .A2(_04922_),
    .B1(_04924_),
    .B2(\as2650.regs[3][2] ),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10048_ (.A1(_02340_),
    .A2(_04920_),
    .B(_04927_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10049_ (.A1(_02387_),
    .A2(_04922_),
    .B1(_04924_),
    .B2(\as2650.regs[3][3] ),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10050_ (.A1(_02386_),
    .A2(_04920_),
    .B(_04928_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10051_ (.I(_04919_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10052_ (.I(_04921_),
    .Z(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10053_ (.I(_04923_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10054_ (.A1(_02432_),
    .A2(_04930_),
    .B1(_04931_),
    .B2(\as2650.regs[3][4] ),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10055_ (.A1(_02431_),
    .A2(_04929_),
    .B(_04932_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10056_ (.A1(_02473_),
    .A2(_04930_),
    .B1(_04931_),
    .B2(\as2650.regs[3][5] ),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10057_ (.A1(_02472_),
    .A2(_04929_),
    .B(_04933_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10058_ (.A1(_02511_),
    .A2(_04930_),
    .B1(_04931_),
    .B2(\as2650.regs[3][6] ),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10059_ (.A1(_02510_),
    .A2(_04929_),
    .B(_04934_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10060_ (.A1(_04757_),
    .A2(_04930_),
    .B1(_04931_),
    .B2(\as2650.regs[3][7] ),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10061_ (.A1(_02553_),
    .A2(_04929_),
    .B(_04935_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10062_ (.A1(_02639_),
    .A2(_02678_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10063_ (.I(_04936_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10064_ (.I(_04937_),
    .Z(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10065_ (.I(_04938_),
    .Z(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10066_ (.I(_04936_),
    .Z(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10067_ (.A1(\as2650.stack[14][0] ),
    .A2(_04940_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10068_ (.A1(_02669_),
    .A2(_04939_),
    .B(_04941_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10069_ (.A1(\as2650.stack[14][1] ),
    .A2(_04940_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10070_ (.A1(_02685_),
    .A2(_04939_),
    .B(_04942_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10071_ (.A1(\as2650.stack[14][2] ),
    .A2(_04940_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10072_ (.A1(_02687_),
    .A2(_04939_),
    .B(_04943_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10073_ (.I(_04937_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10074_ (.A1(\as2650.stack[14][3] ),
    .A2(_04944_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10075_ (.A1(_02689_),
    .A2(_04939_),
    .B(_04945_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10076_ (.I(_04938_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10077_ (.A1(\as2650.stack[14][4] ),
    .A2(_04944_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10078_ (.A1(_02692_),
    .A2(_04946_),
    .B(_04947_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10079_ (.A1(\as2650.stack[14][5] ),
    .A2(_04944_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10080_ (.A1(_02695_),
    .A2(_04946_),
    .B(_04948_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10081_ (.A1(\as2650.stack[14][6] ),
    .A2(_04944_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10082_ (.A1(_02697_),
    .A2(_04946_),
    .B(_04949_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10083_ (.I(_04937_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10084_ (.A1(\as2650.stack[14][7] ),
    .A2(_04950_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10085_ (.A1(_02699_),
    .A2(_04946_),
    .B(_04951_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10086_ (.I(_04937_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10087_ (.A1(\as2650.stack[14][8] ),
    .A2(_04950_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10088_ (.A1(_02702_),
    .A2(_04952_),
    .B(_04953_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10089_ (.A1(\as2650.stack[14][9] ),
    .A2(_04950_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10090_ (.A1(_02705_),
    .A2(_04952_),
    .B(_04954_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10091_ (.A1(\as2650.stack[14][10] ),
    .A2(_04950_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10092_ (.A1(_02707_),
    .A2(_04952_),
    .B(_04955_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10093_ (.A1(\as2650.stack[14][11] ),
    .A2(_04938_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10094_ (.A1(_02709_),
    .A2(_04952_),
    .B(_04956_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10095_ (.A1(\as2650.stack[14][12] ),
    .A2(_04938_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10096_ (.A1(_02711_),
    .A2(_04940_),
    .B(_04957_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10097_ (.A1(_02662_),
    .A2(_02716_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10098_ (.I(_04958_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10099_ (.A1(\as2650.stack[14][13] ),
    .A2(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10100_ (.A1(_02713_),
    .A2(_04959_),
    .B(_04960_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10101_ (.A1(\as2650.stack[14][14] ),
    .A2(_04958_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10102_ (.A1(_02720_),
    .A2(_04959_),
    .B(_04961_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10103_ (.A1(\as2650.stack[14][15] ),
    .A2(_04958_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10104_ (.A1(_02722_),
    .A2(_04959_),
    .B(_04962_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10105_ (.I(_01874_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10106_ (.A1(_01614_),
    .A2(_02558_),
    .A3(_02063_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10107_ (.I(_04964_),
    .Z(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10108_ (.I(_04965_),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10109_ (.I(_04964_),
    .Z(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10110_ (.I(_04967_),
    .Z(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10111_ (.A1(\as2650.stack[13][0] ),
    .A2(_04968_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10112_ (.A1(_04963_),
    .A2(_04966_),
    .B(_04969_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10113_ (.I(_01902_),
    .Z(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10114_ (.A1(\as2650.stack[13][1] ),
    .A2(_04968_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10115_ (.A1(_04970_),
    .A2(_04966_),
    .B(_04971_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10116_ (.I(_01917_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10117_ (.A1(\as2650.stack[13][2] ),
    .A2(_04968_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10118_ (.A1(_04972_),
    .A2(_04966_),
    .B(_04973_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10119_ (.I(_01931_),
    .Z(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10120_ (.A1(\as2650.stack[13][3] ),
    .A2(_04968_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10121_ (.A1(_04974_),
    .A2(_04966_),
    .B(_04975_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10122_ (.I(_01951_),
    .Z(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10123_ (.I(_04965_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10124_ (.I(_04967_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10125_ (.A1(\as2650.stack[13][4] ),
    .A2(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10126_ (.A1(_04976_),
    .A2(_04977_),
    .B(_04979_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10127_ (.I(_01966_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10128_ (.A1(\as2650.stack[13][5] ),
    .A2(_04978_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10129_ (.A1(_04980_),
    .A2(_04977_),
    .B(_04981_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10130_ (.I(_01978_),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10131_ (.A1(\as2650.stack[13][6] ),
    .A2(_04978_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10132_ (.A1(_04982_),
    .A2(_04977_),
    .B(_04983_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10133_ (.I(_01990_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10134_ (.A1(\as2650.stack[13][7] ),
    .A2(_04978_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10135_ (.A1(_04984_),
    .A2(_04977_),
    .B(_04985_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10136_ (.I(_02007_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10137_ (.I(_04965_),
    .Z(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10138_ (.I(_04967_),
    .Z(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(\as2650.stack[13][8] ),
    .A2(_04988_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10140_ (.A1(_04986_),
    .A2(_04987_),
    .B(_04989_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10141_ (.I(_02020_),
    .Z(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10142_ (.A1(\as2650.stack[13][9] ),
    .A2(_04988_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10143_ (.A1(_04990_),
    .A2(_04987_),
    .B(_04991_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10144_ (.I(_02034_),
    .Z(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10145_ (.A1(\as2650.stack[13][10] ),
    .A2(_04988_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10146_ (.A1(_04992_),
    .A2(_04987_),
    .B(_04993_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10147_ (.I(_02047_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10148_ (.A1(\as2650.stack[13][11] ),
    .A2(_04988_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10149_ (.A1(_04994_),
    .A2(_04987_),
    .B(_04995_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10150_ (.I(_02059_),
    .Z(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10151_ (.I(_04965_),
    .Z(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10152_ (.I(_04967_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10153_ (.A1(\as2650.stack[13][12] ),
    .A2(_04998_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10154_ (.A1(_04996_),
    .A2(_04997_),
    .B(_04999_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10155_ (.I(_02070_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10156_ (.A1(\as2650.stack[13][13] ),
    .A2(_04998_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10157_ (.A1(_05000_),
    .A2(_04997_),
    .B(_05001_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10158_ (.I(_02077_),
    .Z(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10159_ (.A1(\as2650.stack[13][14] ),
    .A2(_04998_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10160_ (.A1(_05002_),
    .A2(_04997_),
    .B(_05003_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10161_ (.I(_02084_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10162_ (.A1(\as2650.stack[13][15] ),
    .A2(_04998_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10163_ (.A1(_05004_),
    .A2(_04997_),
    .B(_05005_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10164_ (.A1(_02594_),
    .A2(_02678_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10165_ (.I(_05006_),
    .Z(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10166_ (.I(_05007_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10167_ (.I(_05006_),
    .Z(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10168_ (.I(_05009_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10169_ (.A1(\as2650.stack[12][0] ),
    .A2(_05010_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10170_ (.A1(_04963_),
    .A2(_05008_),
    .B(_05011_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10171_ (.A1(\as2650.stack[12][1] ),
    .A2(_05010_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10172_ (.A1(_04970_),
    .A2(_05008_),
    .B(_05012_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10173_ (.A1(\as2650.stack[12][2] ),
    .A2(_05010_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10174_ (.A1(_04972_),
    .A2(_05008_),
    .B(_05013_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10175_ (.A1(\as2650.stack[12][3] ),
    .A2(_05010_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10176_ (.A1(_04974_),
    .A2(_05008_),
    .B(_05014_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10177_ (.I(_05007_),
    .Z(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10178_ (.I(_05009_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10179_ (.A1(\as2650.stack[12][4] ),
    .A2(_05016_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10180_ (.A1(_04976_),
    .A2(_05015_),
    .B(_05017_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10181_ (.A1(\as2650.stack[12][5] ),
    .A2(_05016_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10182_ (.A1(_04980_),
    .A2(_05015_),
    .B(_05018_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10183_ (.A1(\as2650.stack[12][6] ),
    .A2(_05016_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10184_ (.A1(_04982_),
    .A2(_05015_),
    .B(_05019_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10185_ (.A1(\as2650.stack[12][7] ),
    .A2(_05016_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10186_ (.A1(_04984_),
    .A2(_05015_),
    .B(_05020_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10187_ (.I(_05007_),
    .Z(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10188_ (.I(_05009_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10189_ (.A1(\as2650.stack[12][8] ),
    .A2(_05022_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10190_ (.A1(_04986_),
    .A2(_05021_),
    .B(_05023_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10191_ (.A1(\as2650.stack[12][9] ),
    .A2(_05022_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10192_ (.A1(_04990_),
    .A2(_05021_),
    .B(_05024_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10193_ (.A1(\as2650.stack[12][10] ),
    .A2(_05022_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10194_ (.A1(_04992_),
    .A2(_05021_),
    .B(_05025_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10195_ (.A1(\as2650.stack[12][11] ),
    .A2(_05022_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10196_ (.A1(_04994_),
    .A2(_05021_),
    .B(_05026_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10197_ (.I(_05007_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10198_ (.I(_05009_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10199_ (.A1(\as2650.stack[12][12] ),
    .A2(_05028_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10200_ (.A1(_04996_),
    .A2(_05027_),
    .B(_05029_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10201_ (.A1(\as2650.stack[12][13] ),
    .A2(_05028_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10202_ (.A1(_05000_),
    .A2(_05027_),
    .B(_05030_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10203_ (.A1(\as2650.stack[12][14] ),
    .A2(_05028_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10204_ (.A1(_05002_),
    .A2(_05027_),
    .B(_05031_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10205_ (.A1(\as2650.stack[12][15] ),
    .A2(_05028_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10206_ (.A1(_05004_),
    .A2(_05027_),
    .B(_05032_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10207_ (.A1(_02596_),
    .A2(_04406_),
    .A3(_02595_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10208_ (.A1(_02676_),
    .A2(_05033_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10209_ (.I(_05034_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10210_ (.I(_05035_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10211_ (.I(_05034_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10212_ (.I(_05037_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10213_ (.A1(\as2650.stack[11][0] ),
    .A2(_05038_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10214_ (.A1(_04963_),
    .A2(_05036_),
    .B(_05039_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10215_ (.A1(\as2650.stack[11][1] ),
    .A2(_05038_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10216_ (.A1(_04970_),
    .A2(_05036_),
    .B(_05040_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10217_ (.A1(\as2650.stack[11][2] ),
    .A2(_05038_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10218_ (.A1(_04972_),
    .A2(_05036_),
    .B(_05041_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10219_ (.A1(\as2650.stack[11][3] ),
    .A2(_05038_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10220_ (.A1(_04974_),
    .A2(_05036_),
    .B(_05042_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10221_ (.I(_05035_),
    .Z(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10222_ (.I(_05037_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10223_ (.A1(\as2650.stack[11][4] ),
    .A2(_05044_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10224_ (.A1(_04976_),
    .A2(_05043_),
    .B(_05045_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10225_ (.A1(\as2650.stack[11][5] ),
    .A2(_05044_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10226_ (.A1(_04980_),
    .A2(_05043_),
    .B(_05046_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10227_ (.A1(\as2650.stack[11][6] ),
    .A2(_05044_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10228_ (.A1(_04982_),
    .A2(_05043_),
    .B(_05047_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10229_ (.A1(\as2650.stack[11][7] ),
    .A2(_05044_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10230_ (.A1(_04984_),
    .A2(_05043_),
    .B(_05048_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10231_ (.I(_05035_),
    .Z(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10232_ (.I(_05037_),
    .Z(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10233_ (.A1(\as2650.stack[11][8] ),
    .A2(_05050_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10234_ (.A1(_04986_),
    .A2(_05049_),
    .B(_05051_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10235_ (.A1(\as2650.stack[11][9] ),
    .A2(_05050_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10236_ (.A1(_04990_),
    .A2(_05049_),
    .B(_05052_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10237_ (.A1(\as2650.stack[11][10] ),
    .A2(_05050_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10238_ (.A1(_04992_),
    .A2(_05049_),
    .B(_05053_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10239_ (.A1(\as2650.stack[11][11] ),
    .A2(_05050_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10240_ (.A1(_04994_),
    .A2(_05049_),
    .B(_05054_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10241_ (.I(_05035_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10242_ (.I(_05037_),
    .Z(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10243_ (.A1(\as2650.stack[11][12] ),
    .A2(_05056_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10244_ (.A1(_04996_),
    .A2(_05055_),
    .B(_05057_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10245_ (.I(_02070_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10246_ (.A1(\as2650.stack[11][13] ),
    .A2(_05056_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10247_ (.A1(_05058_),
    .A2(_05055_),
    .B(_05059_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10248_ (.I(_02077_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10249_ (.A1(\as2650.stack[11][14] ),
    .A2(_05056_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10250_ (.A1(_05060_),
    .A2(_05055_),
    .B(_05061_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10251_ (.I(_02084_),
    .Z(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10252_ (.A1(\as2650.stack[11][15] ),
    .A2(_05056_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10253_ (.A1(_05062_),
    .A2(_05055_),
    .B(_05063_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10254_ (.A1(_02179_),
    .A2(_02188_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10255_ (.A1(_04739_),
    .A2(_03913_),
    .A3(_05064_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10256_ (.A1(_04918_),
    .A2(_05065_),
    .B(_02208_),
    .C(_04738_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10257_ (.I(_05066_),
    .Z(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10258_ (.A1(_04918_),
    .A2(_05065_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10259_ (.I(_05068_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10260_ (.A1(_04738_),
    .A2(_02221_),
    .B(_05068_),
    .C(_02222_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10261_ (.I(_05070_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10262_ (.A1(_04841_),
    .A2(_05069_),
    .B1(_05071_),
    .B2(\as2650.regs[6][0] ),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10263_ (.A1(_02170_),
    .A2(_05067_),
    .B(_05072_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10264_ (.A1(_02296_),
    .A2(_05069_),
    .B1(_05071_),
    .B2(\as2650.regs[6][1] ),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10265_ (.A1(_02294_),
    .A2(_05067_),
    .B(_05073_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10266_ (.A1(_02341_),
    .A2(_05069_),
    .B1(_05071_),
    .B2(\as2650.regs[6][2] ),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10267_ (.A1(_02340_),
    .A2(_05067_),
    .B(_05074_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10268_ (.A1(_02387_),
    .A2(_05069_),
    .B1(_05071_),
    .B2(\as2650.regs[6][3] ),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10269_ (.A1(_02386_),
    .A2(_05067_),
    .B(_05075_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10270_ (.I(_05066_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10271_ (.I(_05068_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10272_ (.I(_05070_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10273_ (.A1(_02432_),
    .A2(_05077_),
    .B1(_05078_),
    .B2(\as2650.regs[6][4] ),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10274_ (.A1(_02431_),
    .A2(_05076_),
    .B(_05079_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10275_ (.A1(_02473_),
    .A2(_05077_),
    .B1(_05078_),
    .B2(\as2650.regs[6][5] ),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10276_ (.A1(_02472_),
    .A2(_05076_),
    .B(_05080_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10277_ (.A1(_02511_),
    .A2(_05077_),
    .B1(_05078_),
    .B2(\as2650.regs[6][6] ),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10278_ (.A1(_02510_),
    .A2(_05076_),
    .B(_05081_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10279_ (.A1(_02554_),
    .A2(_05077_),
    .B1(_05078_),
    .B2(\as2650.regs[6][7] ),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10280_ (.A1(_02553_),
    .A2(_05076_),
    .B(_05082_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10281_ (.A1(_02639_),
    .A2(_05033_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10282_ (.I(_05083_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10283_ (.I(_05084_),
    .Z(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10284_ (.I(_05083_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10285_ (.I(_05086_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10286_ (.A1(\as2650.stack[10][0] ),
    .A2(_05087_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10287_ (.A1(_04963_),
    .A2(_05085_),
    .B(_05088_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10288_ (.A1(\as2650.stack[10][1] ),
    .A2(_05087_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10289_ (.A1(_04970_),
    .A2(_05085_),
    .B(_05089_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10290_ (.A1(\as2650.stack[10][2] ),
    .A2(_05087_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10291_ (.A1(_04972_),
    .A2(_05085_),
    .B(_05090_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10292_ (.A1(\as2650.stack[10][3] ),
    .A2(_05087_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10293_ (.A1(_04974_),
    .A2(_05085_),
    .B(_05091_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10294_ (.I(_05084_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10295_ (.I(_05086_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10296_ (.A1(\as2650.stack[10][4] ),
    .A2(_05093_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10297_ (.A1(_04976_),
    .A2(_05092_),
    .B(_05094_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10298_ (.A1(\as2650.stack[10][5] ),
    .A2(_05093_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10299_ (.A1(_04980_),
    .A2(_05092_),
    .B(_05095_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10300_ (.A1(\as2650.stack[10][6] ),
    .A2(_05093_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10301_ (.A1(_04982_),
    .A2(_05092_),
    .B(_05096_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10302_ (.A1(\as2650.stack[10][7] ),
    .A2(_05093_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10303_ (.A1(_04984_),
    .A2(_05092_),
    .B(_05097_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10304_ (.I(_05084_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10305_ (.I(_05086_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10306_ (.A1(\as2650.stack[10][8] ),
    .A2(_05099_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10307_ (.A1(_04986_),
    .A2(_05098_),
    .B(_05100_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10308_ (.A1(\as2650.stack[10][9] ),
    .A2(_05099_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10309_ (.A1(_04990_),
    .A2(_05098_),
    .B(_05101_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10310_ (.A1(\as2650.stack[10][10] ),
    .A2(_05099_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10311_ (.A1(_04992_),
    .A2(_05098_),
    .B(_05102_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10312_ (.A1(\as2650.stack[10][11] ),
    .A2(_05099_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10313_ (.A1(_04994_),
    .A2(_05098_),
    .B(_05103_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10314_ (.I(_05084_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10315_ (.I(_05086_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10316_ (.A1(\as2650.stack[10][12] ),
    .A2(_05105_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10317_ (.A1(_04996_),
    .A2(_05104_),
    .B(_05106_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10318_ (.A1(\as2650.stack[10][13] ),
    .A2(_05105_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10319_ (.A1(_05058_),
    .A2(_05104_),
    .B(_05107_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10320_ (.A1(\as2650.stack[10][14] ),
    .A2(_05105_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10321_ (.A1(_05060_),
    .A2(_05104_),
    .B(_05108_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10322_ (.A1(\as2650.stack[10][15] ),
    .A2(_05105_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10323_ (.A1(_05062_),
    .A2(_05104_),
    .B(_05109_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10324_ (.I(_01874_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10325_ (.A1(_01876_),
    .A2(_01883_),
    .A3(_03149_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10326_ (.I(_05111_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10327_ (.I(_05112_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10328_ (.I(_05113_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10329_ (.I(_05111_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10330_ (.A1(\as2650.stack[0][0] ),
    .A2(_05115_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10331_ (.A1(_05110_),
    .A2(_05114_),
    .B(_05116_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10332_ (.I(_01902_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10333_ (.A1(\as2650.stack[0][1] ),
    .A2(_05115_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10334_ (.A1(_05117_),
    .A2(_05114_),
    .B(_05118_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10335_ (.I(_01917_),
    .Z(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10336_ (.A1(\as2650.stack[0][2] ),
    .A2(_05115_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10337_ (.A1(_05119_),
    .A2(_05114_),
    .B(_05120_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10338_ (.I(_01931_),
    .Z(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10339_ (.I(_05112_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10340_ (.A1(\as2650.stack[0][3] ),
    .A2(_05122_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10341_ (.A1(_05121_),
    .A2(_05114_),
    .B(_05123_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10342_ (.I(_01951_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10343_ (.I(_05113_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10344_ (.A1(\as2650.stack[0][4] ),
    .A2(_05122_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10345_ (.A1(_05124_),
    .A2(_05125_),
    .B(_05126_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10346_ (.I(_01966_),
    .Z(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10347_ (.A1(\as2650.stack[0][5] ),
    .A2(_05122_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10348_ (.A1(_05127_),
    .A2(_05125_),
    .B(_05128_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10349_ (.I(_01978_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10350_ (.A1(\as2650.stack[0][6] ),
    .A2(_05122_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10351_ (.A1(_05129_),
    .A2(_05125_),
    .B(_05130_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10352_ (.I(_01990_),
    .Z(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10353_ (.I(_05112_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10354_ (.A1(\as2650.stack[0][7] ),
    .A2(_05132_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10355_ (.A1(_05131_),
    .A2(_05125_),
    .B(_05133_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10356_ (.I(_02007_),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10357_ (.I(_05112_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10358_ (.A1(\as2650.stack[0][8] ),
    .A2(_05132_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10359_ (.A1(_05134_),
    .A2(_05135_),
    .B(_05136_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10360_ (.I(_02020_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10361_ (.A1(\as2650.stack[0][9] ),
    .A2(_05132_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10362_ (.A1(_05137_),
    .A2(_05135_),
    .B(_05138_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10363_ (.I(_02034_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10364_ (.A1(\as2650.stack[0][10] ),
    .A2(_05132_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10365_ (.A1(_05139_),
    .A2(_05135_),
    .B(_05140_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10366_ (.I(_02047_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10367_ (.A1(\as2650.stack[0][11] ),
    .A2(_05113_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10368_ (.A1(_05141_),
    .A2(_05135_),
    .B(_05142_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10369_ (.I(_02059_),
    .Z(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10370_ (.A1(\as2650.stack[0][12] ),
    .A2(_05113_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10371_ (.A1(_05143_),
    .A2(_05115_),
    .B(_05144_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10372_ (.A1(_02595_),
    .A2(_03132_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10373_ (.I(_05145_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10374_ (.A1(\as2650.stack[0][13] ),
    .A2(_05146_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10375_ (.A1(_05000_),
    .A2(_05146_),
    .B(_05147_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10376_ (.A1(\as2650.stack[0][14] ),
    .A2(_05145_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10377_ (.A1(_05002_),
    .A2(_05146_),
    .B(_05148_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10378_ (.A1(\as2650.stack[0][15] ),
    .A2(_05145_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10379_ (.A1(_05004_),
    .A2(_05146_),
    .B(_05149_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10380_ (.A1(_02594_),
    .A2(_05033_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10381_ (.I(_05150_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10382_ (.I(_05151_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10383_ (.I(_05150_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10384_ (.I(_05153_),
    .Z(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(\as2650.stack[8][0] ),
    .A2(_05154_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10386_ (.A1(_05110_),
    .A2(_05152_),
    .B(_05155_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10387_ (.A1(\as2650.stack[8][1] ),
    .A2(_05154_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10388_ (.A1(_05117_),
    .A2(_05152_),
    .B(_05156_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10389_ (.A1(\as2650.stack[8][2] ),
    .A2(_05154_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10390_ (.A1(_05119_),
    .A2(_05152_),
    .B(_05157_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10391_ (.A1(\as2650.stack[8][3] ),
    .A2(_05154_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10392_ (.A1(_05121_),
    .A2(_05152_),
    .B(_05158_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10393_ (.I(_05151_),
    .Z(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10394_ (.I(_05153_),
    .Z(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10395_ (.A1(\as2650.stack[8][4] ),
    .A2(_05160_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10396_ (.A1(_05124_),
    .A2(_05159_),
    .B(_05161_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10397_ (.A1(\as2650.stack[8][5] ),
    .A2(_05160_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10398_ (.A1(_05127_),
    .A2(_05159_),
    .B(_05162_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10399_ (.A1(\as2650.stack[8][6] ),
    .A2(_05160_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10400_ (.A1(_05129_),
    .A2(_05159_),
    .B(_05163_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10401_ (.A1(\as2650.stack[8][7] ),
    .A2(_05160_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10402_ (.A1(_05131_),
    .A2(_05159_),
    .B(_05164_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10403_ (.I(_05151_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10404_ (.I(_05153_),
    .Z(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10405_ (.A1(\as2650.stack[8][8] ),
    .A2(_05166_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10406_ (.A1(_05134_),
    .A2(_05165_),
    .B(_05167_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10407_ (.A1(\as2650.stack[8][9] ),
    .A2(_05166_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10408_ (.A1(_05137_),
    .A2(_05165_),
    .B(_05168_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10409_ (.A1(\as2650.stack[8][10] ),
    .A2(_05166_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10410_ (.A1(_05139_),
    .A2(_05165_),
    .B(_05169_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10411_ (.A1(\as2650.stack[8][11] ),
    .A2(_05166_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10412_ (.A1(_05141_),
    .A2(_05165_),
    .B(_05170_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10413_ (.I(_05151_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10414_ (.I(_05153_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10415_ (.A1(\as2650.stack[8][12] ),
    .A2(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10416_ (.A1(_05143_),
    .A2(_05171_),
    .B(_05173_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10417_ (.A1(\as2650.stack[8][13] ),
    .A2(_05172_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10418_ (.A1(_05058_),
    .A2(_05171_),
    .B(_05174_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10419_ (.A1(\as2650.stack[8][14] ),
    .A2(_05172_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10420_ (.A1(_05060_),
    .A2(_05171_),
    .B(_05175_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10421_ (.A1(\as2650.stack[8][15] ),
    .A2(_05172_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10422_ (.A1(_05062_),
    .A2(_05171_),
    .B(_05176_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10423_ (.A1(_02599_),
    .A2(_02676_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10424_ (.I(_05177_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10425_ (.I(_05178_),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10426_ (.I(_05179_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10427_ (.I(_05177_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10428_ (.A1(\as2650.stack[7][0] ),
    .A2(_05181_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10429_ (.A1(_05110_),
    .A2(_05180_),
    .B(_05182_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10430_ (.A1(\as2650.stack[7][1] ),
    .A2(_05181_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10431_ (.A1(_05117_),
    .A2(_05180_),
    .B(_05183_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10432_ (.A1(\as2650.stack[7][2] ),
    .A2(_05181_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10433_ (.A1(_05119_),
    .A2(_05180_),
    .B(_05184_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10434_ (.I(_05178_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10435_ (.A1(\as2650.stack[7][3] ),
    .A2(_05185_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10436_ (.A1(_05121_),
    .A2(_05180_),
    .B(_05186_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10437_ (.I(_05179_),
    .Z(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10438_ (.A1(\as2650.stack[7][4] ),
    .A2(_05185_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10439_ (.A1(_05124_),
    .A2(_05187_),
    .B(_05188_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10440_ (.A1(\as2650.stack[7][5] ),
    .A2(_05185_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10441_ (.A1(_05127_),
    .A2(_05187_),
    .B(_05189_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10442_ (.A1(\as2650.stack[7][6] ),
    .A2(_05185_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10443_ (.A1(_05129_),
    .A2(_05187_),
    .B(_05190_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10444_ (.I(_05178_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10445_ (.A1(\as2650.stack[7][7] ),
    .A2(_05191_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10446_ (.A1(_05131_),
    .A2(_05187_),
    .B(_05192_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10447_ (.I(_05178_),
    .Z(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10448_ (.A1(\as2650.stack[7][8] ),
    .A2(_05191_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10449_ (.A1(_05134_),
    .A2(_05193_),
    .B(_05194_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10450_ (.A1(\as2650.stack[7][9] ),
    .A2(_05191_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10451_ (.A1(_05137_),
    .A2(_05193_),
    .B(_05195_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10452_ (.A1(\as2650.stack[7][10] ),
    .A2(_05191_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10453_ (.A1(_05139_),
    .A2(_05193_),
    .B(_05196_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10454_ (.A1(\as2650.stack[7][11] ),
    .A2(_05179_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10455_ (.A1(_05141_),
    .A2(_05193_),
    .B(_05197_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10456_ (.A1(\as2650.stack[7][12] ),
    .A2(_05179_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10457_ (.A1(_05143_),
    .A2(_05181_),
    .B(_05198_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10458_ (.A1(_02627_),
    .A2(_02715_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10459_ (.I(_05199_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10460_ (.A1(\as2650.stack[7][13] ),
    .A2(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10461_ (.A1(_05000_),
    .A2(_05200_),
    .B(_05201_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10462_ (.A1(\as2650.stack[7][14] ),
    .A2(_05199_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10463_ (.A1(_05002_),
    .A2(_05200_),
    .B(_05202_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10464_ (.A1(\as2650.stack[7][15] ),
    .A2(_05199_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10465_ (.A1(_05004_),
    .A2(_05200_),
    .B(_05203_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10466_ (.A1(_02557_),
    .A2(_02558_),
    .A3(_02063_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10467_ (.I(_05204_),
    .Z(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10468_ (.I(_05205_),
    .Z(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10469_ (.I(_05204_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10470_ (.I(_05207_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10471_ (.A1(\as2650.stack[9][0] ),
    .A2(_05208_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10472_ (.A1(_05110_),
    .A2(_05206_),
    .B(_05209_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10473_ (.A1(\as2650.stack[9][1] ),
    .A2(_05208_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10474_ (.A1(_05117_),
    .A2(_05206_),
    .B(_05210_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10475_ (.A1(\as2650.stack[9][2] ),
    .A2(_05208_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10476_ (.A1(_05119_),
    .A2(_05206_),
    .B(_05211_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10477_ (.A1(\as2650.stack[9][3] ),
    .A2(_05208_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10478_ (.A1(_05121_),
    .A2(_05206_),
    .B(_05212_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10479_ (.I(_05205_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10480_ (.I(_05207_),
    .Z(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10481_ (.A1(\as2650.stack[9][4] ),
    .A2(_05214_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10482_ (.A1(_05124_),
    .A2(_05213_),
    .B(_05215_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10483_ (.A1(\as2650.stack[9][5] ),
    .A2(_05214_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10484_ (.A1(_05127_),
    .A2(_05213_),
    .B(_05216_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10485_ (.A1(\as2650.stack[9][6] ),
    .A2(_05214_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10486_ (.A1(_05129_),
    .A2(_05213_),
    .B(_05217_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10487_ (.A1(\as2650.stack[9][7] ),
    .A2(_05214_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10488_ (.A1(_05131_),
    .A2(_05213_),
    .B(_05218_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10489_ (.I(_05205_),
    .Z(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10490_ (.I(_05207_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10491_ (.A1(\as2650.stack[9][8] ),
    .A2(_05220_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10492_ (.A1(_05134_),
    .A2(_05219_),
    .B(_05221_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10493_ (.A1(\as2650.stack[9][9] ),
    .A2(_05220_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10494_ (.A1(_05137_),
    .A2(_05219_),
    .B(_05222_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10495_ (.A1(\as2650.stack[9][10] ),
    .A2(_05220_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10496_ (.A1(_05139_),
    .A2(_05219_),
    .B(_05223_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10497_ (.A1(\as2650.stack[9][11] ),
    .A2(_05220_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10498_ (.A1(_05141_),
    .A2(_05219_),
    .B(_05224_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10499_ (.I(_05205_),
    .Z(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10500_ (.I(_05207_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10501_ (.A1(\as2650.stack[9][12] ),
    .A2(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10502_ (.A1(_05143_),
    .A2(_05225_),
    .B(_05227_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10503_ (.A1(\as2650.stack[9][13] ),
    .A2(_05226_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10504_ (.A1(_05058_),
    .A2(_05225_),
    .B(_05228_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10505_ (.A1(\as2650.stack[9][14] ),
    .A2(_05226_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10506_ (.A1(_05060_),
    .A2(_05225_),
    .B(_05229_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10507_ (.A1(\as2650.stack[9][15] ),
    .A2(_05226_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10508_ (.A1(_05062_),
    .A2(_05225_),
    .B(_05230_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10509_ (.D(_00011_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10510_ (.D(_00012_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(net106));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10511_ (.D(_00013_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(net107));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10512_ (.D(_00014_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(net118));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10513_ (.D(_00015_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(net129));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10514_ (.D(_00016_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10515_ (.D(_00017_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10516_ (.D(_00018_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10517_ (.D(_00019_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10518_ (.D(_00020_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10519_ (.D(_00021_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10520_ (.D(_00022_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(net138));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10521_ (.D(_00023_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(net108));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10522_ (.D(_00024_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net109));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10523_ (.D(_00025_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net110));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10524_ (.D(_00026_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net111));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10525_ (.D(_00027_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net112));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10526_ (.D(_00028_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(net113));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10527_ (.D(_00029_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(net114));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10528_ (.D(_00030_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(net115));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10529_ (.D(_00031_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(net116));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10530_ (.D(_00032_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(net117));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10531_ (.D(_00033_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(net119));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10532_ (.D(_00034_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(net120));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10533_ (.D(_00035_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(net121));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10534_ (.D(_00036_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(net122));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10535_ (.D(_00037_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(net123));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10536_ (.D(_00038_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(net124));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10537_ (.D(_00039_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(net125));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10538_ (.D(_00040_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(net126));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10539_ (.D(_00041_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(net127));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10540_ (.D(_00042_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(net128));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10541_ (.D(_00043_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(net130));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10542_ (.D(_00044_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(net131));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10543_ (.D(_00045_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10544_ (.D(net343),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10545_ (.D(net377),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(wb_debug_carry));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10546_ (.D(net332),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\web_behavior[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10547_ (.D(net309),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\web_behavior[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10548_ (.D(_00050_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\wb_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10549_ (.D(net367),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\wb_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10550_ (.D(_00052_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\wb_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10551_ (.D(_00053_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\wb_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10552_ (.D(net306),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\wb_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10553_ (.D(net274),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\wb_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10554_ (.D(net270),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\wb_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10555_ (.D(net266),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\wb_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10556_ (.D(net286),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\wb_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10557_ (.D(net340),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\wb_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10558_ (.D(net290),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\wb_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10559_ (.D(net278),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\wb_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10560_ (.D(net282),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\wb_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10561_ (.D(net373),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\wb_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10562_ (.D(net364),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\wb_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10563_ (.D(net349),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\wb_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10564_ (.D(net358),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\wb_counter[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10565_ (.D(_00067_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\wb_counter[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10566_ (.D(net370),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\wb_counter[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10567_ (.D(net346),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\wb_counter[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10568_ (.D(net355),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\wb_counter[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10569_ (.D(net361),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\wb_counter[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10570_ (.D(net352),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\wb_counter[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10571_ (.D(net298),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\wb_counter[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10572_ (.D(net325),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\wb_counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10573_ (.D(net321),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\wb_counter[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10574_ (.D(net313),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\wb_counter[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10575_ (.D(net302),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\wb_counter[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10576_ (.D(net317),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\wb_counter[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10577_ (.D(net329),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\wb_counter[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10578_ (.D(net294),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\wb_counter[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10579_ (.D(net336),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\wb_counter[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10580_ (.D(_00082_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10581_ (.D(_00083_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10582_ (.D(_00084_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10583_ (.D(_00085_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10584_ (.D(_00086_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10585_ (.D(_00087_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10586_ (.D(_00088_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10587_ (.D(_00089_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10588_ (.D(_00090_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10589_ (.D(_00091_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10590_ (.D(_00092_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10591_ (.D(_00093_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10592_ (.D(_00094_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10593_ (.D(_00095_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10594_ (.D(_00096_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10595_ (.D(_00097_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10596_ (.D(_00098_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10597_ (.D(_00099_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10598_ (.D(_00100_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10599_ (.D(_00101_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10600_ (.D(_00102_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.regs[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10601_ (.D(_00103_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.regs[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10602_ (.D(_00104_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10603_ (.D(_00105_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10604_ (.D(_00106_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10605_ (.D(_00107_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10606_ (.D(_00108_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10607_ (.D(_00109_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10608_ (.D(_00110_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10609_ (.D(_00111_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10610_ (.D(_00112_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10611_ (.D(_00113_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10612_ (.D(_00114_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10613_ (.D(_00115_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10614_ (.D(_00116_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10615_ (.D(_00117_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10616_ (.D(_00118_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10617_ (.D(_00119_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10618_ (.D(_00120_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10619_ (.D(_00121_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10620_ (.D(_00122_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10621_ (.D(_00123_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10622_ (.D(_00124_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10623_ (.D(_00125_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10624_ (.D(_00126_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10625_ (.D(_00127_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10626_ (.D(_00128_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10627_ (.D(_00129_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10628_ (.D(_00130_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10629_ (.D(_00131_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10630_ (.D(_00132_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10631_ (.D(_00133_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10632_ (.D(_00134_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10633_ (.D(_00135_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10634_ (.D(_00136_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10635_ (.D(_00137_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10636_ (.D(_00138_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10637_ (.D(_00139_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10638_ (.D(_00140_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10639_ (.D(_00141_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10640_ (.D(_00142_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10641_ (.D(_00143_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10642_ (.D(_00144_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10643_ (.D(_00145_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10644_ (.D(_00146_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10645_ (.D(_00147_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10646_ (.D(_00148_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10647_ (.D(_00149_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10648_ (.D(_00150_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10649_ (.D(_00151_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10650_ (.D(_00152_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10651_ (.D(_00153_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10652_ (.D(_00154_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10653_ (.D(_00155_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10654_ (.D(_00156_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10655_ (.D(_00157_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10656_ (.D(_00158_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10657_ (.D(_00159_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10658_ (.D(_00160_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10659_ (.D(_00161_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10660_ (.D(_00162_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10661_ (.D(_00163_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10662_ (.D(_00164_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10663_ (.D(_00165_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10664_ (.D(_00166_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10665_ (.D(_00167_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10666_ (.D(_00168_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10667_ (.D(_00169_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10668_ (.D(_00170_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10669_ (.D(_00171_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10670_ (.D(_00172_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10671_ (.D(_00173_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10672_ (.D(_00174_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10673_ (.D(_00175_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10674_ (.D(_00176_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10675_ (.D(_00177_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10676_ (.D(_00178_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10677_ (.D(_00179_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10678_ (.D(_00180_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10679_ (.D(_00181_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10680_ (.D(_00182_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10681_ (.D(_00183_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10682_ (.D(_00184_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10683_ (.D(_00185_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _10684_ (.D(_00007_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10685_ (.D(_00005_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10686_ (.D(_00008_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10687_ (.D(_00009_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10688_ (.D(_00006_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10689_ (.D(net139),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10690_ (.D(_00186_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.last_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10691_ (.D(_00187_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.last_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10692_ (.D(_00188_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.last_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10693_ (.D(_00189_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.last_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10694_ (.D(_00190_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.last_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10695_ (.D(_00191_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.last_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10696_ (.D(_00192_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.last_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10697_ (.D(_00193_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.last_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10698_ (.D(_00194_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10699_ (.D(_00195_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10700_ (.D(_00196_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10701_ (.D(_00197_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10702_ (.D(_00198_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10703_ (.D(_00199_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10704_ (.D(_00200_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10705_ (.D(_00201_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10706_ (.D(_00202_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10707_ (.D(_00203_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10708_ (.D(_00204_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10709_ (.D(_00205_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10710_ (.D(_00206_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10711_ (.D(_00207_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10712_ (.D(_00208_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10713_ (.D(_00209_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10714_ (.D(_00210_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.chirp_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10715_ (.D(_00211_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.chirp_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10716_ (.D(_00212_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.chirp_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10717_ (.D(_00213_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.indirect_target[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10718_ (.D(_00214_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.indirect_target[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10719_ (.D(_00215_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.indirect_target[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10720_ (.D(_00216_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.indirect_target[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10721_ (.D(_00217_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\as2650.indirect_target[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10722_ (.D(_00218_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.indirect_target[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10723_ (.D(_00219_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.indirect_target[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10724_ (.D(_00220_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.indirect_target[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10725_ (.D(_00221_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.indirect_target[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10726_ (.D(_00222_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.indirect_target[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10727_ (.D(_00223_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.indirect_target[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10728_ (.D(_00224_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.indirect_target[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10729_ (.D(_00225_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.indirect_target[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10730_ (.D(_00226_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10731_ (.D(_00227_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10732_ (.D(_00228_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10733_ (.D(_00229_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.indexed_cyc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10734_ (.D(_00230_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(\as2650.indexed_cyc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10735_ (.D(_00231_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.indirect_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10736_ (.D(_00232_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.extend ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10737_ (.D(_00233_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(net98));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10738_ (.D(_00234_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10739_ (.D(_00235_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10740_ (.D(_00236_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.instruction_args_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10741_ (.D(_00237_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10742_ (.D(_00238_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.instruction_args_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10743_ (.D(_00239_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10744_ (.D(_00240_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10745_ (.D(_00241_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.instruction_args_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10746_ (.D(_00242_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10747_ (.D(_00243_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10748_ (.D(_00244_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10749_ (.D(_00245_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10750_ (.D(_00246_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10751_ (.D(_00247_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10752_ (.D(_00248_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10753_ (.D(_00249_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.instruction_args_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10754_ (.D(_00250_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.instruction_args_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10755_ (.D(_00251_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10756_ (.D(_00252_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10757_ (.D(_00253_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10758_ (.D(_00254_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10759_ (.D(_00255_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.insin[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10760_ (.D(_00256_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.insin[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10761_ (.D(_00257_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.insin[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10762_ (.D(_00258_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.insin[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10763_ (.D(_00259_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.insin[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10764_ (.D(_00260_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.insin[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10765_ (.D(_00261_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10766_ (.D(_00262_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.insin[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10767_ (.D(_00263_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.last_addr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10768_ (.D(_00264_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.last_addr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10769_ (.D(_00265_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.last_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10770_ (.D(_00266_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.last_addr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10771_ (.D(_00267_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.last_addr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10772_ (.D(_00268_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.last_addr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10773_ (.D(_00269_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.last_addr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10774_ (.D(_00270_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.last_addr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10775_ (.D(_00271_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.PC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10776_ (.D(_00272_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10777_ (.D(_00273_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10778_ (.D(_00274_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.PC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10779_ (.D(_00275_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10780_ (.D(_00276_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10781_ (.D(_00277_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10782_ (.D(_00278_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10783_ (.D(_00279_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10784_ (.D(_00280_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10785_ (.D(_00281_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10786_ (.D(_00282_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10787_ (.D(_00283_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10788_ (.D(_00284_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.debug_psl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10789_ (.D(_00285_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10790_ (.D(_00286_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10791_ (.D(_00287_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10792_ (.D(_00288_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10793_ (.D(_00289_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.debug_psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10794_ (.D(_00290_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.debug_psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10795_ (.D(_00291_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10796_ (.D(_00292_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.debug_psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10797_ (.D(_00293_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.debug_psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10798_ (.D(_00294_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.debug_psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10799_ (.D(_00295_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10800_ (.D(_00296_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10801_ (.D(_00297_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10802_ (.D(_00298_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10803_ (.D(_00299_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10804_ (.D(_00300_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.chirpchar[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10805_ (.D(_00301_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.regs[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10806_ (.D(_00302_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\as2650.regs[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10807_ (.D(_00303_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.regs[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10808_ (.D(_00304_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10809_ (.D(_00305_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10810_ (.D(_00306_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10811_ (.D(_00307_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10812_ (.D(_00308_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10813_ (.D(_00309_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10814_ (.D(_00310_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10815_ (.D(_00311_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.regs[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10816_ (.D(_00312_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10817_ (.D(_00313_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.regs[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10818_ (.D(_00314_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.regs[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10819_ (.D(_00315_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10820_ (.D(_00316_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10821_ (.D(_00317_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.chirpchar[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10822_ (.D(_00000_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.chirpchar[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10823_ (.D(_00001_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.chirpchar[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10824_ (.D(_00002_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.chirpchar[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10825_ (.D(_00003_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.chirpchar[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10826_ (.D(_00004_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.chirpchar[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10827_ (.D(_00318_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10828_ (.D(_00319_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10829_ (.D(_00320_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10830_ (.D(_00321_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10831_ (.D(_00322_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10832_ (.D(_00323_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.regs[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10833_ (.D(_00324_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10834_ (.D(_00325_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10835_ (.D(_00326_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10836_ (.D(_00327_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10837_ (.D(_00328_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10838_ (.D(_00329_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10839_ (.D(_00330_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10840_ (.D(_00331_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10841_ (.D(_00332_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10842_ (.D(_00333_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10843_ (.D(_00334_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10844_ (.D(_00335_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10845_ (.D(_00336_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10846_ (.D(_00337_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10847_ (.D(_00338_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10848_ (.D(_00339_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10849_ (.D(_00340_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10850_ (.D(_00341_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10851_ (.D(_00342_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\as2650.regs[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10852_ (.D(_00343_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10853_ (.D(_00344_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10854_ (.D(_00345_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10855_ (.D(_00346_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10856_ (.D(_00347_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _10857_ (.D(_00348_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10858_ (.D(_00349_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.regs[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10859_ (.D(_00350_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10860_ (.D(_00351_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10861_ (.D(_00352_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10862_ (.D(_00353_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10863_ (.D(_00354_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10864_ (.D(_00355_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10865_ (.D(_00356_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10866_ (.D(_00357_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10867_ (.D(_00358_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10868_ (.D(_00359_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10869_ (.D(_00360_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10870_ (.D(_00361_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10871_ (.D(_00362_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10872_ (.D(_00363_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10873_ (.D(_00364_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10874_ (.D(_00365_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10875_ (.D(_00366_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10876_ (.D(_00367_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10877_ (.D(_00368_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10878_ (.D(_00369_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10879_ (.D(_00370_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10880_ (.D(_00371_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10881_ (.D(_00372_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10882_ (.D(_00373_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10883_ (.D(_00374_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10884_ (.D(_00375_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10885_ (.D(_00376_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10886_ (.D(_00377_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10887_ (.D(_00378_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10888_ (.D(_00379_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10889_ (.D(_00380_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10890_ (.D(_00381_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10891_ (.D(_00382_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10892_ (.D(_00383_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10893_ (.D(_00384_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10894_ (.D(_00385_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10895_ (.D(_00386_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10896_ (.D(_00387_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10897_ (.D(_00388_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10898_ (.D(_00389_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10899_ (.D(_00390_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10900_ (.D(_00391_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10901_ (.D(_00392_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10902_ (.D(_00393_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10903_ (.D(_00394_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10904_ (.D(_00395_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10905_ (.D(_00396_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10906_ (.D(_00397_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10907_ (.D(_00398_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10908_ (.D(_00399_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10909_ (.D(_00400_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10910_ (.D(_00401_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10911_ (.D(_00402_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10912_ (.D(_00403_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10913_ (.D(_00404_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10914_ (.D(_00405_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10915_ (.D(_00406_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10916_ (.D(_00407_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10917_ (.D(_00408_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10918_ (.D(_00409_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10919_ (.D(_00410_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10920_ (.D(_00411_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10921_ (.D(_00412_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10922_ (.D(_00413_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10923_ (.D(_00414_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10924_ (.D(_00415_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10925_ (.D(_00416_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10926_ (.D(_00417_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10927_ (.D(_00418_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.regs[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10928_ (.D(_00419_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.regs[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10929_ (.D(_00420_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.regs[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10930_ (.D(_00421_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10931_ (.D(_00422_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10932_ (.D(_00423_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10933_ (.D(_00424_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10934_ (.D(_00425_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10935_ (.D(_00426_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10936_ (.D(_00427_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10937_ (.D(_00428_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10938_ (.D(_00429_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10939_ (.D(_00430_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10940_ (.D(_00431_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10941_ (.D(_00432_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10942_ (.D(_00433_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10943_ (.D(_00434_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10944_ (.D(_00435_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10945_ (.D(_00436_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10946_ (.D(_00437_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10947_ (.D(_00438_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10948_ (.D(_00439_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10949_ (.D(_00440_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10950_ (.D(_00441_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10951_ (.D(_00442_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10952_ (.D(_00443_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10953_ (.D(_00444_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10954_ (.D(_00445_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10955_ (.D(_00446_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10956_ (.D(_00447_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10957_ (.D(_00448_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10958_ (.D(_00449_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10959_ (.D(_00450_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10960_ (.D(_00451_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10961_ (.D(_00452_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10962_ (.D(_00453_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10963_ (.D(_00454_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10964_ (.D(_00455_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10965_ (.D(_00456_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10966_ (.D(_00457_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10967_ (.D(_00458_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10968_ (.D(_00459_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10969_ (.D(_00460_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10970_ (.D(_00461_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10971_ (.D(_00462_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10972_ (.D(_00463_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10973_ (.D(_00464_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10974_ (.D(_00465_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10975_ (.D(_00466_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10976_ (.D(_00467_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10977_ (.D(_00468_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10978_ (.D(_00469_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10979_ (.D(_00470_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10980_ (.D(_00471_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10981_ (.D(_00472_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10982_ (.D(_00473_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10983_ (.D(_00474_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10984_ (.D(_00475_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10985_ (.D(_00476_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10986_ (.D(_00477_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10987_ (.D(_00478_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10988_ (.D(_00479_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10989_ (.D(_00480_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10990_ (.D(_00481_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10991_ (.D(_00482_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10992_ (.D(_00483_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10993_ (.D(_00484_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10994_ (.D(_00485_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10995_ (.D(_00486_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10996_ (.D(_00487_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10997_ (.D(_00488_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10998_ (.D(_00489_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10999_ (.D(_00490_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11000_ (.D(_00491_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11001_ (.D(_00492_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11002_ (.D(_00493_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11003_ (.D(_00494_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11004_ (.D(_00495_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11005_ (.D(_00496_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11006_ (.D(_00497_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11007_ (.D(_00498_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11008_ (.D(_00499_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11009_ (.D(_00500_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11010_ (.D(_00501_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11097_ (.I(net141),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11098_ (.I(net141),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11099_ (.I(net141),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11100_ (.I(net142),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11101_ (.I(net142),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11102_ (.I(net142),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11103_ (.I(net143),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11104_ (.I(net141),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0__01311_ (.I(_01311_),
    .Z(clknet_0__01311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f__01311_ (.I(clknet_0__01311_),
    .Z(clknet_1_0__leaf__01311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f__01311_ (.I(clknet_0__01311_),
    .Z(clknet_1_1__leaf__01311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_110_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_118_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_128_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_129_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_84_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_90_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout142 (.I(net51),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout143 (.I(net51),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout144 (.I(net67),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold100 (.I(_01705_),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(_00048_),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(wbs_dat_i[31]),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold103 (.I(net39),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold104 (.I(_01839_),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold105 (.I(_00081_),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold106 (.I(wbs_dat_i[9]),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold107 (.I(net46),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold108 (.I(_01753_),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold109 (.I(_00059_),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold110 (.I(net389),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold111 (.I(_01700_),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold112 (.I(_00046_),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold113 (.I(wbs_dat_i[19]),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold114 (.I(_01792_),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold115 (.I(_00069_),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold116 (.I(wbs_dat_i[15]),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold117 (.I(_01775_),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold118 (.I(_00065_),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold119 (.I(wbs_dat_i[22]),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold120 (.I(_01805_),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold121 (.I(_00072_),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold122 (.I(wbs_dat_i[20]),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold123 (.I(_01796_),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold124 (.I(_00070_),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold125 (.I(wbs_dat_i[16]),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold126 (.I(_01778_),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold127 (.I(_00066_),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold128 (.I(wbs_dat_i[21]),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold129 (.I(_01802_),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold130 (.I(_00071_),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold131 (.I(wbs_dat_i[14]),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold132 (.I(_01772_),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold133 (.I(_00064_),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold134 (.I(wbs_dat_i[1]),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold135 (.I(_01717_),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold136 (.I(_00051_),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold137 (.I(wbs_dat_i[18]),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold138 (.I(_01789_),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold139 (.I(_00068_),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold140 (.I(wbs_dat_i[13]),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold141 (.I(_01768_),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold142 (.I(_00063_),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold143 (.I(wbs_adr_i[22]),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold144 (.I(wbs_adr_i[21]),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold145 (.I(_01697_),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold146 (.I(_00047_),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold147 (.I(net387),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold148 (.I(wbs_cyc_i),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold149 (.I(_01557_),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold150 (.I(wbs_dat_i[17]),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold151 (.I(wbs_dat_i[2]),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold152 (.I(wbs_dat_i[0]),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold153 (.I(wbs_dat_i[3]),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold154 (.I(_01724_),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(wbs_dat_i[7]),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(net44),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(_01742_),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(_00057_),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(wbs_dat_i[6]),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(net43),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(_01739_),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(_00056_),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(wbs_dat_i[5]),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(net42),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(_01736_),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(_00055_),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(wbs_dat_i[11]),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(net17),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(_01759_),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(_00061_),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(wbs_dat_i[12]),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(net18),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(_01762_),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(_00062_),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(wbs_dat_i[8]),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(net45),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(_01746_),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(_00058_),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(wbs_dat_i[10]),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(net16),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(_01757_),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(_00060_),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(wbs_dat_i[30]),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(net38),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(_01836_),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(_00080_),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(wbs_dat_i[23]),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(net30),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(_01809_),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(_00073_),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(wbs_dat_i[27]),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(net34),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(_01825_),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(_00077_),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(wbs_dat_i[4]),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(net41),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(_01728_),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(_00054_),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(net390),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(_01707_),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(_00049_),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(wbs_dat_i[26]),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(net33),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(_01822_),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(_00076_),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(wbs_dat_i[28]),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(net35),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(_01828_),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(_00078_),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(wbs_dat_i[25]),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(net32),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(_01818_),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(_00075_),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(wbs_dat_i[24]),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(net31),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(_01812_),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(_00074_),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(wbs_dat_i[29]),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(net36),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(_01833_),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold98 (.I(_00079_),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(net388),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(io_in[9]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(wb_rst_i),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(net375),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input13 (.I(net374),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(net379),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input15 (.I(net341),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(net287),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(net275),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(net279),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(net371),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input2 (.I(io_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(net362),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(net347),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(net356),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(net378),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(net368),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(net344),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input26 (.I(net365),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(net353),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(net359),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(net350),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(io_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(net295),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(net322),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(net318),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(net310),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(net299),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(net314),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(net326),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input37 (.I(net330),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(net291),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(net333),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(io_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input40 (.I(net307),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(net303),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(net271),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(net267),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(net263),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(net283),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input46 (.I(net337),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(wbs_stb_i),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(wbs_we_i),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(io_in[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input6 (.I(io_in[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input7 (.I(io_in[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input8 (.I(io_in[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input9 (.I(io_in[8]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output100 (.I(net100),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output101 (.I(net101),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output102 (.I(net102),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output103 (.I(net103),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output104 (.I(net104),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output105 (.I(net105),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output124 (.I(net124),
    .Z(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output125 (.I(net125),
    .Z(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output126 (.I(net126),
    .Z(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output127 (.I(net127),
    .Z(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output128 (.I(net128),
    .Z(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output129 (.I(net129),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output130 (.I(net130),
    .Z(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output131 (.I(net131),
    .Z(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output132 (.I(net132),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output133 (.I(net133),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output134 (.I(net134),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output135 (.I(net135),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output136 (.I(net136),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output137 (.I(net137),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output138 (.I(net138),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output49 (.I(net49),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output50 (.I(net50),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output51 (.I(net143),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output52 (.I(net52),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output53 (.I(net53),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output54 (.I(net54),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output55 (.I(net55),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output56 (.I(net56),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output57 (.I(net57),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output58 (.I(net58),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output59 (.I(net59),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output60 (.I(net60),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output61 (.I(net61),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output62 (.I(net62),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output63 (.I(net63),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output64 (.I(net64),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output65 (.I(net65),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output66 (.I(net66),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output67 (.I(net144),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output68 (.I(net68),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output69 (.I(net69),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output70 (.I(net70),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output71 (.I(net71),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output72 (.I(net72),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output73 (.I(net73),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output74 (.I(net74),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output75 (.I(net75),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output76 (.I(net76),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output77 (.I(net77),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output78 (.I(net78),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output79 (.I(net79),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output80 (.I(net80),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output81 (.I(net81),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output82 (.I(net82),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output83 (.I(net83),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output84 (.I(net84),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output85 (.I(net85),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output86 (.I(net86),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output87 (.I(net87),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output88 (.I(net88),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output89 (.I(net89),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output90 (.I(net90),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output91 (.I(net91),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output92 (.I(net92),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output93 (.I(net93),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output94 (.I(net94),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output95 (.I(net95),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output96 (.I(net96),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output97 (.I(net97),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output98 (.I(net98),
    .Z(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output99 (.I(net99),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer1 (.I(net236),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 rebuffer10 (.I(_00913_),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer11 (.I(_00638_),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer12 (.I(_00873_),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer13 (.I(net243),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer14 (.I(net254),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer15 (.I(net245),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer16 (.I(net246),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer17 (.I(_00708_),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer18 (.I(_00811_),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer19 (.I(_00907_),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer2 (.I(net232),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer20 (.I(_01238_),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer21 (.I(_02968_),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer22 (.I(_00892_),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer23 (.I(net256),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer24 (.I(_00823_),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer25 (.I(_00701_),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer26 (.I(_00842_),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer27 (.I(_00989_),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer28 (.I(_00700_),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer29 (.I(_00757_),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer3 (.I(net383),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer30 (.I(_00897_),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer31 (.I(_00719_),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer32 (.I(_01169_),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer33 (.I(_00875_),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer34 (.I(_00719_),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer35 (.I(_00860_),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer36 (.I(_00658_),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer37 (.I(_01246_),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer4 (.I(_00818_),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_00981_),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer6 (.I(_00887_),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer7 (.I(_00783_),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer8 (.I(net242),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer9 (.I(_00638_),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire139 (.I(net140),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire140 (.I(_00010_),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_194 (.Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_195 (.Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_196 (.Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_197 (.Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_198 (.Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_199 (.Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_200 (.Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_201 (.Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_202 (.Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_203 (.Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_204 (.Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_205 (.Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_206 (.Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_207 (.Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_208 (.Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_209 (.Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_210 (.Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_211 (.Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_212 (.Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_213 (.Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_214 (.Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_215 (.Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_216 (.Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_217 (.Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_218 (.Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_219 (.Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_220 (.Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_221 (.Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_222 (.Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_223 (.Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_224 (.Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_225 (.Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_226 (.Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_227 (.Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_228 (.Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_229 (.Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_230 (.Z(net230));
 assign io_oeb[0] = net194;
 assign io_oeb[13] = net147;
 assign io_oeb[14] = net148;
 assign io_oeb[15] = net149;
 assign io_oeb[16] = net150;
 assign io_oeb[17] = net151;
 assign io_oeb[18] = net152;
 assign io_oeb[19] = net197;
 assign io_oeb[1] = net145;
 assign io_oeb[20] = net198;
 assign io_oeb[21] = net199;
 assign io_oeb[22] = net200;
 assign io_oeb[23] = net201;
 assign io_oeb[24] = net202;
 assign io_oeb[25] = net203;
 assign io_oeb[26] = net204;
 assign io_oeb[27] = net205;
 assign io_oeb[28] = net206;
 assign io_oeb[29] = net207;
 assign io_oeb[2] = net146;
 assign io_oeb[30] = net208;
 assign io_oeb[31] = net209;
 assign io_oeb[32] = net210;
 assign io_oeb[33] = net211;
 assign io_oeb[34] = net212;
 assign io_oeb[35] = net213;
 assign io_oeb[36] = net214;
 assign io_oeb[37] = net215;
 assign io_oeb[3] = net195;
 assign io_oeb[4] = net196;
 assign io_out[0] = net153;
 assign io_out[19] = net156;
 assign io_out[20] = net157;
 assign io_out[21] = net158;
 assign io_out[22] = net159;
 assign io_out[23] = net160;
 assign io_out[24] = net161;
 assign io_out[25] = net162;
 assign io_out[26] = net163;
 assign io_out[27] = net164;
 assign io_out[28] = net165;
 assign io_out[29] = net166;
 assign io_out[30] = net167;
 assign io_out[31] = net168;
 assign io_out[32] = net169;
 assign io_out[33] = net170;
 assign io_out[34] = net171;
 assign io_out[35] = net172;
 assign io_out[36] = net173;
 assign io_out[37] = net174;
 assign io_out[3] = net154;
 assign io_out[4] = net155;
 assign irq[0] = net175;
 assign irq[1] = net176;
 assign irq[2] = net177;
 assign la_data_out[33] = net178;
 assign la_data_out[34] = net179;
 assign la_data_out[35] = net180;
 assign la_data_out[36] = net181;
 assign la_data_out[37] = net182;
 assign la_data_out[38] = net183;
 assign la_data_out[39] = net184;
 assign la_data_out[40] = net185;
 assign la_data_out[41] = net216;
 assign la_data_out[42] = net217;
 assign la_data_out[43] = net218;
 assign la_data_out[44] = net219;
 assign la_data_out[45] = net220;
 assign la_data_out[46] = net221;
 assign la_data_out[47] = net222;
 assign la_data_out[48] = net223;
 assign la_data_out[49] = net186;
 assign la_data_out[50] = net187;
 assign la_data_out[51] = net188;
 assign la_data_out[52] = net189;
 assign la_data_out[53] = net190;
 assign la_data_out[54] = net191;
 assign la_data_out[55] = net192;
 assign la_data_out[56] = net193;
 assign la_data_out[57] = net224;
 assign la_data_out[58] = net225;
 assign la_data_out[59] = net226;
 assign la_data_out[60] = net227;
 assign la_data_out[61] = net228;
 assign la_data_out[62] = net229;
 assign la_data_out[63] = net230;
endmodule

