magic
tech gf180mcuD
magscale 1 10
timestamp 1701963987
<< metal1 >>
rect 20178 46398 20190 46450
rect 20242 46447 20254 46450
rect 20962 46447 20974 46450
rect 20242 46401 20974 46447
rect 20242 46398 20254 46401
rect 20962 46398 20974 46401
rect 21026 46398 21038 46450
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 26238 46114 26290 46126
rect 26238 46050 26290 46062
rect 29486 46114 29538 46126
rect 29486 46050 29538 46062
rect 33182 46114 33234 46126
rect 33182 46050 33234 46062
rect 36990 46114 37042 46126
rect 36990 46050 37042 46062
rect 40798 46114 40850 46126
rect 40798 46050 40850 46062
rect 44606 46114 44658 46126
rect 44606 46050 44658 46062
rect 1934 46002 1986 46014
rect 1934 45938 1986 45950
rect 6638 46002 6690 46014
rect 6638 45938 6690 45950
rect 7198 46002 7250 46014
rect 7198 45938 7250 45950
rect 8094 46002 8146 46014
rect 8094 45938 8146 45950
rect 10782 46002 10834 46014
rect 10782 45938 10834 45950
rect 13470 46002 13522 46014
rect 13470 45938 13522 45950
rect 14814 46002 14866 46014
rect 14814 45938 14866 45950
rect 16382 46002 16434 46014
rect 16382 45938 16434 45950
rect 18846 46002 18898 46014
rect 18846 45938 18898 45950
rect 20190 46002 20242 46014
rect 20190 45938 20242 45950
rect 22878 46002 22930 46014
rect 22878 45938 22930 45950
rect 47630 46002 47682 46014
rect 47630 45938 47682 45950
rect 5630 45890 5682 45902
rect 4274 45838 4286 45890
rect 4338 45838 4350 45890
rect 4722 45838 4734 45890
rect 4786 45838 4798 45890
rect 5630 45826 5682 45838
rect 6190 45890 6242 45902
rect 6190 45826 6242 45838
rect 9662 45890 9714 45902
rect 9662 45826 9714 45838
rect 11006 45890 11058 45902
rect 11006 45826 11058 45838
rect 12238 45890 12290 45902
rect 12238 45826 12290 45838
rect 13694 45890 13746 45902
rect 13694 45826 13746 45838
rect 15038 45890 15090 45902
rect 17726 45890 17778 45902
rect 48190 45890 48242 45902
rect 17042 45838 17054 45890
rect 17106 45838 17118 45890
rect 19282 45838 19294 45890
rect 19346 45838 19358 45890
rect 20962 45838 20974 45890
rect 21026 45838 21038 45890
rect 21970 45838 21982 45890
rect 22034 45838 22046 45890
rect 23314 45838 23326 45890
rect 23378 45838 23390 45890
rect 25218 45838 25230 45890
rect 25282 45838 25294 45890
rect 28914 45838 28926 45890
rect 28978 45838 28990 45890
rect 32162 45838 32174 45890
rect 32226 45838 32238 45890
rect 35970 45838 35982 45890
rect 36034 45838 36046 45890
rect 39778 45838 39790 45890
rect 39842 45838 39854 45890
rect 43922 45838 43934 45890
rect 43986 45838 43998 45890
rect 15038 45826 15090 45838
rect 17726 45826 17778 45838
rect 48190 45826 48242 45838
rect 8766 45778 8818 45790
rect 8766 45714 8818 45726
rect 4958 45666 5010 45678
rect 4958 45602 5010 45614
rect 8430 45666 8482 45678
rect 8430 45602 8482 45614
rect 9998 45666 10050 45678
rect 9998 45602 10050 45614
rect 11342 45666 11394 45678
rect 15374 45666 15426 45678
rect 18062 45666 18114 45678
rect 12562 45614 12574 45666
rect 12626 45614 12638 45666
rect 14018 45614 14030 45666
rect 14082 45614 14094 45666
rect 17266 45614 17278 45666
rect 17330 45614 17342 45666
rect 11342 45602 11394 45614
rect 15374 45602 15426 45614
rect 18062 45602 18114 45614
rect 19070 45666 19122 45678
rect 19070 45602 19122 45614
rect 20750 45666 20802 45678
rect 20750 45602 20802 45614
rect 21758 45666 21810 45678
rect 21758 45602 21810 45614
rect 23102 45666 23154 45678
rect 23102 45602 23154 45614
rect 47854 45666 47906 45678
rect 47854 45602 47906 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 9662 45330 9714 45342
rect 12798 45330 12850 45342
rect 11666 45278 11678 45330
rect 11730 45278 11742 45330
rect 9662 45266 9714 45278
rect 12798 45266 12850 45278
rect 17614 45330 17666 45342
rect 17614 45266 17666 45278
rect 21534 45330 21586 45342
rect 21534 45266 21586 45278
rect 28142 45330 28194 45342
rect 28142 45266 28194 45278
rect 31838 45330 31890 45342
rect 31838 45266 31890 45278
rect 36990 45330 37042 45342
rect 36990 45266 37042 45278
rect 41918 45330 41970 45342
rect 41918 45266 41970 45278
rect 44830 45330 44882 45342
rect 44830 45266 44882 45278
rect 7534 45218 7586 45230
rect 7534 45154 7586 45166
rect 7870 45218 7922 45230
rect 7870 45154 7922 45166
rect 8654 45218 8706 45230
rect 8654 45154 8706 45166
rect 25902 45218 25954 45230
rect 25902 45154 25954 45166
rect 12014 45106 12066 45118
rect 3938 45054 3950 45106
rect 4002 45054 4014 45106
rect 7186 45054 7198 45106
rect 7250 45054 7262 45106
rect 8418 45054 8430 45106
rect 8482 45054 8494 45106
rect 12014 45042 12066 45054
rect 25566 45106 25618 45118
rect 27122 45054 27134 45106
rect 27186 45054 27198 45106
rect 31602 45054 31614 45106
rect 31666 45054 31678 45106
rect 35186 45054 35198 45106
rect 35250 45054 35262 45106
rect 35970 45054 35982 45106
rect 36034 45054 36046 45106
rect 41010 45054 41022 45106
rect 41074 45054 41086 45106
rect 43810 45054 43822 45106
rect 43874 45054 43886 45106
rect 25566 45042 25618 45054
rect 4846 44994 4898 45006
rect 4846 44930 4898 44942
rect 30158 44994 30210 45006
rect 30158 44930 30210 44942
rect 33294 44994 33346 45006
rect 33294 44930 33346 44942
rect 1934 44882 1986 44894
rect 1934 44818 1986 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 25454 44546 25506 44558
rect 30830 44546 30882 44558
rect 28466 44494 28478 44546
rect 28530 44494 28542 44546
rect 25454 44482 25506 44494
rect 30830 44482 30882 44494
rect 37998 44546 38050 44558
rect 37998 44482 38050 44494
rect 40910 44546 40962 44558
rect 40910 44482 40962 44494
rect 45838 44546 45890 44558
rect 45838 44482 45890 44494
rect 15262 44434 15314 44446
rect 27470 44434 27522 44446
rect 1922 44382 1934 44434
rect 1986 44382 1998 44434
rect 8866 44382 8878 44434
rect 8930 44382 8942 44434
rect 16370 44382 16382 44434
rect 16434 44382 16446 44434
rect 27906 44382 27918 44434
rect 27970 44382 27982 44434
rect 15262 44370 15314 44382
rect 27470 44370 27522 44382
rect 14702 44322 14754 44334
rect 28254 44322 28306 44334
rect 4834 44270 4846 44322
rect 4898 44270 4910 44322
rect 5954 44270 5966 44322
rect 6018 44270 6030 44322
rect 19170 44270 19182 44322
rect 19234 44270 19246 44322
rect 24434 44270 24446 44322
rect 24498 44270 24510 44322
rect 29362 44270 29374 44322
rect 29426 44270 29438 44322
rect 29922 44270 29934 44322
rect 29986 44270 29998 44322
rect 35410 44270 35422 44322
rect 35474 44270 35486 44322
rect 36978 44270 36990 44322
rect 37042 44270 37054 44322
rect 39890 44270 39902 44322
rect 39954 44270 39966 44322
rect 44818 44270 44830 44322
rect 44882 44270 44894 44322
rect 14702 44258 14754 44270
rect 28254 44258 28306 44270
rect 22430 44210 22482 44222
rect 4050 44158 4062 44210
rect 4114 44158 4126 44210
rect 6738 44158 6750 44210
rect 6802 44158 6814 44210
rect 11330 44158 11342 44210
rect 11394 44158 11406 44210
rect 18498 44158 18510 44210
rect 18562 44158 18574 44210
rect 22430 44146 22482 44158
rect 22766 44210 22818 44222
rect 22766 44146 22818 44158
rect 23774 44210 23826 44222
rect 23774 44146 23826 44158
rect 24110 44210 24162 44222
rect 24110 44146 24162 44158
rect 29150 44210 29202 44222
rect 29150 44146 29202 44158
rect 32734 44210 32786 44222
rect 32734 44146 32786 44158
rect 33070 44210 33122 44222
rect 33070 44146 33122 44158
rect 33406 44210 33458 44222
rect 33406 44146 33458 44158
rect 33742 44210 33794 44222
rect 33742 44146 33794 44158
rect 34078 44210 34130 44222
rect 34078 44146 34130 44158
rect 34414 44210 34466 44222
rect 34414 44146 34466 44158
rect 35646 44210 35698 44222
rect 35646 44146 35698 44158
rect 42814 44210 42866 44222
rect 42814 44146 42866 44158
rect 43150 44210 43202 44222
rect 43150 44146 43202 44158
rect 43486 44210 43538 44222
rect 43486 44146 43538 44158
rect 43822 44210 43874 44222
rect 43822 44146 43874 44158
rect 9326 44098 9378 44110
rect 9326 44034 9378 44046
rect 11678 44098 11730 44110
rect 11678 44034 11730 44046
rect 14814 44098 14866 44110
rect 14814 44034 14866 44046
rect 15150 44098 15202 44110
rect 15150 44034 15202 44046
rect 19742 44098 19794 44110
rect 19742 44034 19794 44046
rect 21534 44098 21586 44110
rect 21534 44034 21586 44046
rect 21870 44098 21922 44110
rect 21870 44034 21922 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 5294 43762 5346 43774
rect 5294 43698 5346 43710
rect 29934 43762 29986 43774
rect 29934 43698 29986 43710
rect 6750 43650 6802 43662
rect 6750 43586 6802 43598
rect 7422 43650 7474 43662
rect 7422 43586 7474 43598
rect 8094 43650 8146 43662
rect 8094 43586 8146 43598
rect 10558 43650 10610 43662
rect 10558 43586 10610 43598
rect 17950 43650 18002 43662
rect 33406 43650 33458 43662
rect 20962 43598 20974 43650
rect 21026 43598 21038 43650
rect 31602 43598 31614 43650
rect 31666 43598 31678 43650
rect 17950 43586 18002 43598
rect 33406 43586 33458 43598
rect 45278 43650 45330 43662
rect 45278 43586 45330 43598
rect 4734 43538 4786 43550
rect 7870 43538 7922 43550
rect 4274 43486 4286 43538
rect 4338 43486 4350 43538
rect 6962 43486 6974 43538
rect 7026 43486 7038 43538
rect 4734 43474 4786 43486
rect 7870 43474 7922 43486
rect 8206 43538 8258 43550
rect 8206 43474 8258 43486
rect 10446 43538 10498 43550
rect 18062 43538 18114 43550
rect 31278 43538 31330 43550
rect 44942 43538 44994 43550
rect 11330 43486 11342 43538
rect 11394 43486 11406 43538
rect 21298 43486 21310 43538
rect 21362 43486 21374 43538
rect 25330 43486 25342 43538
rect 25394 43486 25406 43538
rect 29586 43486 29598 43538
rect 29650 43486 29662 43538
rect 30146 43486 30158 43538
rect 30210 43486 30222 43538
rect 33170 43486 33182 43538
rect 33234 43486 33246 43538
rect 45602 43486 45614 43538
rect 45666 43486 45678 43538
rect 10446 43474 10498 43486
rect 18062 43474 18114 43486
rect 31278 43474 31330 43486
rect 44942 43474 44994 43486
rect 5630 43426 5682 43438
rect 14814 43426 14866 43438
rect 12114 43374 12126 43426
rect 12178 43374 12190 43426
rect 14242 43374 14254 43426
rect 14306 43374 14318 43426
rect 5630 43362 5682 43374
rect 14814 43362 14866 43374
rect 18510 43426 18562 43438
rect 18510 43362 18562 43374
rect 19182 43426 19234 43438
rect 19182 43362 19234 43374
rect 20414 43426 20466 43438
rect 28702 43426 28754 43438
rect 22082 43374 22094 43426
rect 22146 43374 22158 43426
rect 24210 43374 24222 43426
rect 24274 43374 24286 43426
rect 26002 43374 26014 43426
rect 26066 43374 26078 43426
rect 28130 43374 28142 43426
rect 28194 43374 28206 43426
rect 20414 43362 20466 43374
rect 28702 43362 28754 43374
rect 29038 43426 29090 43438
rect 29038 43362 29090 43374
rect 44606 43426 44658 43438
rect 44606 43362 44658 43374
rect 46622 43426 46674 43438
rect 46622 43362 46674 43374
rect 1934 43314 1986 43326
rect 1934 43250 1986 43262
rect 7534 43314 7586 43326
rect 7534 43250 7586 43262
rect 10558 43314 10610 43326
rect 10558 43250 10610 43262
rect 17950 43314 18002 43326
rect 17950 43250 18002 43262
rect 19406 43314 19458 43326
rect 20638 43314 20690 43326
rect 19730 43262 19742 43314
rect 19794 43262 19806 43314
rect 19406 43250 19458 43262
rect 20638 43250 20690 43262
rect 29262 43314 29314 43326
rect 29262 43250 29314 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 23998 42978 24050 42990
rect 41582 42978 41634 42990
rect 24322 42926 24334 42978
rect 24386 42926 24398 42978
rect 23998 42914 24050 42926
rect 41582 42914 41634 42926
rect 41918 42978 41970 42990
rect 47058 42926 47070 42978
rect 47122 42926 47134 42978
rect 41918 42914 41970 42926
rect 18398 42866 18450 42878
rect 2034 42814 2046 42866
rect 2098 42814 2110 42866
rect 12674 42814 12686 42866
rect 12738 42814 12750 42866
rect 15026 42814 15038 42866
rect 15090 42814 15102 42866
rect 18398 42802 18450 42814
rect 21422 42866 21474 42878
rect 21422 42802 21474 42814
rect 22542 42866 22594 42878
rect 22542 42802 22594 42814
rect 24782 42866 24834 42878
rect 24782 42802 24834 42814
rect 8766 42754 8818 42766
rect 18174 42754 18226 42766
rect 4274 42702 4286 42754
rect 4338 42702 4350 42754
rect 4722 42702 4734 42754
rect 4786 42702 4798 42754
rect 9874 42702 9886 42754
rect 9938 42702 9950 42754
rect 17826 42702 17838 42754
rect 17890 42702 17902 42754
rect 8766 42690 8818 42702
rect 18174 42690 18226 42702
rect 22094 42754 22146 42766
rect 22094 42690 22146 42702
rect 22318 42754 22370 42766
rect 22318 42690 22370 42702
rect 22878 42754 22930 42766
rect 22878 42690 22930 42702
rect 23774 42754 23826 42766
rect 23774 42690 23826 42702
rect 28478 42754 28530 42766
rect 40898 42702 40910 42754
rect 40962 42702 40974 42754
rect 45602 42702 45614 42754
rect 45666 42702 45678 42754
rect 28478 42690 28530 42702
rect 7758 42642 7810 42654
rect 7758 42578 7810 42590
rect 8094 42642 8146 42654
rect 13582 42642 13634 42654
rect 18622 42642 18674 42654
rect 10546 42590 10558 42642
rect 10610 42590 10622 42642
rect 17154 42590 17166 42642
rect 17218 42590 17230 42642
rect 8094 42578 8146 42590
rect 13582 42578 13634 42590
rect 18622 42578 18674 42590
rect 18846 42642 18898 42654
rect 18846 42578 18898 42590
rect 21758 42642 21810 42654
rect 21758 42578 21810 42590
rect 21870 42642 21922 42654
rect 21870 42578 21922 42590
rect 22766 42642 22818 42654
rect 22766 42578 22818 42590
rect 39790 42642 39842 42654
rect 40786 42590 40798 42642
rect 40850 42590 40862 42642
rect 39790 42578 39842 42590
rect 4958 42530 5010 42542
rect 4958 42466 5010 42478
rect 8430 42530 8482 42542
rect 8430 42466 8482 42478
rect 8654 42530 8706 42542
rect 8654 42466 8706 42478
rect 9326 42530 9378 42542
rect 9326 42466 9378 42478
rect 19406 42530 19458 42542
rect 19406 42466 19458 42478
rect 19966 42530 20018 42542
rect 19966 42466 20018 42478
rect 23438 42530 23490 42542
rect 23438 42466 23490 42478
rect 29262 42530 29314 42542
rect 29262 42466 29314 42478
rect 40238 42530 40290 42542
rect 40238 42466 40290 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 10558 42194 10610 42206
rect 10558 42130 10610 42142
rect 11790 42194 11842 42206
rect 11790 42130 11842 42142
rect 17726 42194 17778 42206
rect 17726 42130 17778 42142
rect 22318 42194 22370 42206
rect 22318 42130 22370 42142
rect 7870 42082 7922 42094
rect 7870 42018 7922 42030
rect 8430 42082 8482 42094
rect 8430 42018 8482 42030
rect 8878 42082 8930 42094
rect 8878 42018 8930 42030
rect 9886 42082 9938 42094
rect 9886 42018 9938 42030
rect 9998 42082 10050 42094
rect 9998 42018 10050 42030
rect 10222 42082 10274 42094
rect 10222 42018 10274 42030
rect 18174 42082 18226 42094
rect 18174 42018 18226 42030
rect 18398 42082 18450 42094
rect 18398 42018 18450 42030
rect 18510 42082 18562 42094
rect 18510 42018 18562 42030
rect 22206 42082 22258 42094
rect 22206 42018 22258 42030
rect 7086 41970 7138 41982
rect 3826 41918 3838 41970
rect 3890 41918 3902 41970
rect 7086 41906 7138 41918
rect 7310 41970 7362 41982
rect 7310 41906 7362 41918
rect 7646 41970 7698 41982
rect 7646 41906 7698 41918
rect 7982 41970 8034 41982
rect 7982 41906 8034 41918
rect 8206 41970 8258 41982
rect 8206 41906 8258 41918
rect 8654 41970 8706 41982
rect 8654 41906 8706 41918
rect 8990 41970 9042 41982
rect 8990 41906 9042 41918
rect 10334 41970 10386 41982
rect 10334 41906 10386 41918
rect 10782 41970 10834 41982
rect 10782 41906 10834 41918
rect 10894 41970 10946 41982
rect 10894 41906 10946 41918
rect 11342 41970 11394 41982
rect 11342 41906 11394 41918
rect 11678 41970 11730 41982
rect 11678 41906 11730 41918
rect 11902 41970 11954 41982
rect 11902 41906 11954 41918
rect 16942 41970 16994 41982
rect 16942 41906 16994 41918
rect 17390 41970 17442 41982
rect 17390 41906 17442 41918
rect 17726 41970 17778 41982
rect 17726 41906 17778 41918
rect 18062 41970 18114 41982
rect 18062 41906 18114 41918
rect 22542 41970 22594 41982
rect 22542 41906 22594 41918
rect 23214 41970 23266 41982
rect 23214 41906 23266 41918
rect 23438 41970 23490 41982
rect 23438 41906 23490 41918
rect 23550 41970 23602 41982
rect 23550 41906 23602 41918
rect 23886 41970 23938 41982
rect 27906 41918 27918 41970
rect 27970 41918 27982 41970
rect 23886 41906 23938 41918
rect 7422 41858 7474 41870
rect 4498 41806 4510 41858
rect 4562 41806 4574 41858
rect 6626 41806 6638 41858
rect 6690 41806 6702 41858
rect 7422 41794 7474 41806
rect 22878 41858 22930 41870
rect 31166 41858 31218 41870
rect 28578 41806 28590 41858
rect 28642 41806 28654 41858
rect 30706 41806 30718 41858
rect 30770 41806 30782 41858
rect 22878 41794 22930 41806
rect 31166 41794 31218 41806
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 11902 41410 11954 41422
rect 11902 41346 11954 41358
rect 12462 41410 12514 41422
rect 12462 41346 12514 41358
rect 18622 41410 18674 41422
rect 18622 41346 18674 41358
rect 23214 41410 23266 41422
rect 23214 41346 23266 41358
rect 9214 41298 9266 41310
rect 4834 41246 4846 41298
rect 4898 41246 4910 41298
rect 9214 41234 9266 41246
rect 23774 41298 23826 41310
rect 23774 41234 23826 41246
rect 28030 41298 28082 41310
rect 28030 41234 28082 41246
rect 12014 41186 12066 41198
rect 2034 41134 2046 41186
rect 2098 41134 2110 41186
rect 8306 41134 8318 41186
rect 8370 41134 8382 41186
rect 12014 41122 12066 41134
rect 12574 41186 12626 41198
rect 12574 41122 12626 41134
rect 17838 41186 17890 41198
rect 22878 41186 22930 41198
rect 20290 41134 20302 41186
rect 20354 41134 20366 41186
rect 17838 41122 17890 41134
rect 22878 41122 22930 41134
rect 27582 41186 27634 41198
rect 27582 41122 27634 41134
rect 28254 41186 28306 41198
rect 28254 41122 28306 41134
rect 11566 41074 11618 41086
rect 2706 41022 2718 41074
rect 2770 41022 2782 41074
rect 8082 41022 8094 41074
rect 8146 41022 8158 41074
rect 11566 41010 11618 41022
rect 11902 41074 11954 41086
rect 11902 41010 11954 41022
rect 18174 41074 18226 41086
rect 18174 41010 18226 41022
rect 18734 41074 18786 41086
rect 22542 41074 22594 41086
rect 20066 41022 20078 41074
rect 20130 41022 20142 41074
rect 18734 41010 18786 41022
rect 22542 41010 22594 41022
rect 23102 41074 23154 41086
rect 23102 41010 23154 41022
rect 27806 41074 27858 41086
rect 27806 41010 27858 41022
rect 47630 41074 47682 41086
rect 47630 41010 47682 41022
rect 48190 41074 48242 41086
rect 48190 41010 48242 41022
rect 5742 40962 5794 40974
rect 5742 40898 5794 40910
rect 6862 40962 6914 40974
rect 6862 40898 6914 40910
rect 12462 40962 12514 40974
rect 12462 40898 12514 40910
rect 13694 40962 13746 40974
rect 13694 40898 13746 40910
rect 17726 40962 17778 40974
rect 17726 40898 17778 40910
rect 18062 40962 18114 40974
rect 18062 40898 18114 40910
rect 18622 40962 18674 40974
rect 18622 40898 18674 40910
rect 19294 40962 19346 40974
rect 19294 40898 19346 40910
rect 22318 40962 22370 40974
rect 22318 40898 22370 40910
rect 22654 40962 22706 40974
rect 22654 40898 22706 40910
rect 23214 40962 23266 40974
rect 23214 40898 23266 40910
rect 28590 40962 28642 40974
rect 28590 40898 28642 40910
rect 47854 40962 47906 40974
rect 47854 40898 47906 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 8990 40626 9042 40638
rect 13582 40626 13634 40638
rect 13010 40574 13022 40626
rect 13074 40574 13086 40626
rect 8990 40562 9042 40574
rect 13582 40562 13634 40574
rect 13806 40626 13858 40638
rect 13806 40562 13858 40574
rect 14366 40626 14418 40638
rect 26574 40626 26626 40638
rect 20402 40574 20414 40626
rect 20466 40574 20478 40626
rect 14366 40562 14418 40574
rect 26574 40562 26626 40574
rect 27806 40626 27858 40638
rect 27806 40562 27858 40574
rect 28142 40626 28194 40638
rect 28142 40562 28194 40574
rect 28366 40626 28418 40638
rect 28366 40562 28418 40574
rect 29150 40626 29202 40638
rect 29150 40562 29202 40574
rect 6750 40514 6802 40526
rect 6750 40450 6802 40462
rect 7086 40514 7138 40526
rect 7086 40450 7138 40462
rect 8430 40514 8482 40526
rect 8430 40450 8482 40462
rect 8542 40514 8594 40526
rect 8542 40450 8594 40462
rect 27022 40514 27074 40526
rect 27022 40450 27074 40462
rect 27582 40514 27634 40526
rect 27582 40450 27634 40462
rect 8206 40402 8258 40414
rect 4274 40350 4286 40402
rect 4338 40350 4350 40402
rect 8206 40338 8258 40350
rect 13358 40402 13410 40414
rect 13358 40338 13410 40350
rect 13918 40402 13970 40414
rect 26910 40402 26962 40414
rect 20626 40350 20638 40402
rect 20690 40350 20702 40402
rect 13918 40338 13970 40350
rect 26910 40338 26962 40350
rect 27246 40402 27298 40414
rect 27246 40338 27298 40350
rect 27470 40402 27522 40414
rect 27470 40338 27522 40350
rect 28030 40402 28082 40414
rect 28030 40338 28082 40350
rect 28814 40402 28866 40414
rect 28814 40338 28866 40350
rect 32510 40290 32562 40302
rect 32510 40226 32562 40238
rect 1934 40178 1986 40190
rect 1934 40114 1986 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 15038 39730 15090 39742
rect 15038 39666 15090 39678
rect 15374 39730 15426 39742
rect 15374 39666 15426 39678
rect 15710 39730 15762 39742
rect 15710 39666 15762 39678
rect 16830 39730 16882 39742
rect 16830 39666 16882 39678
rect 26126 39730 26178 39742
rect 26126 39666 26178 39678
rect 28142 39730 28194 39742
rect 30146 39678 30158 39730
rect 30210 39678 30222 39730
rect 32274 39678 32286 39730
rect 32338 39678 32350 39730
rect 35522 39678 35534 39730
rect 35586 39678 35598 39730
rect 28142 39666 28194 39678
rect 7086 39618 7138 39630
rect 7086 39554 7138 39566
rect 7310 39618 7362 39630
rect 7310 39554 7362 39566
rect 14590 39618 14642 39630
rect 14590 39554 14642 39566
rect 23326 39618 23378 39630
rect 23326 39554 23378 39566
rect 27246 39618 27298 39630
rect 27246 39554 27298 39566
rect 27582 39618 27634 39630
rect 27582 39554 27634 39566
rect 27918 39618 27970 39630
rect 27918 39554 27970 39566
rect 28254 39618 28306 39630
rect 28254 39554 28306 39566
rect 28478 39618 28530 39630
rect 35982 39618 36034 39630
rect 29474 39566 29486 39618
rect 29538 39566 29550 39618
rect 32722 39566 32734 39618
rect 32786 39566 32798 39618
rect 39554 39566 39566 39618
rect 39618 39566 39630 39618
rect 28478 39554 28530 39566
rect 35982 39554 36034 39566
rect 6750 39506 6802 39518
rect 6750 39442 6802 39454
rect 14702 39506 14754 39518
rect 14702 39442 14754 39454
rect 21982 39506 22034 39518
rect 23774 39506 23826 39518
rect 22306 39454 22318 39506
rect 22370 39454 22382 39506
rect 21982 39442 22034 39454
rect 23774 39442 23826 39454
rect 23998 39506 24050 39518
rect 23998 39442 24050 39454
rect 26462 39506 26514 39518
rect 26462 39442 26514 39454
rect 26574 39506 26626 39518
rect 33394 39454 33406 39506
rect 33458 39454 33470 39506
rect 26574 39442 26626 39454
rect 6974 39394 7026 39406
rect 6974 39330 7026 39342
rect 14142 39394 14194 39406
rect 14142 39330 14194 39342
rect 14254 39394 14306 39406
rect 14254 39330 14306 39342
rect 14814 39394 14866 39406
rect 14814 39330 14866 39342
rect 16270 39394 16322 39406
rect 16270 39330 16322 39342
rect 17390 39394 17442 39406
rect 17390 39330 17442 39342
rect 17838 39394 17890 39406
rect 17838 39330 17890 39342
rect 21310 39394 21362 39406
rect 23662 39394 23714 39406
rect 21634 39342 21646 39394
rect 21698 39342 21710 39394
rect 21310 39330 21362 39342
rect 23662 39330 23714 39342
rect 26798 39394 26850 39406
rect 26798 39330 26850 39342
rect 27358 39394 27410 39406
rect 39778 39342 39790 39394
rect 39842 39342 39854 39394
rect 27358 39330 27410 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 10222 39058 10274 39070
rect 10222 38994 10274 39006
rect 12014 39058 12066 39070
rect 12014 38994 12066 39006
rect 12574 39058 12626 39070
rect 12574 38994 12626 39006
rect 13918 39058 13970 39070
rect 13918 38994 13970 39006
rect 14478 39058 14530 39070
rect 25342 39058 25394 39070
rect 16818 39006 16830 39058
rect 16882 39006 16894 39058
rect 14478 38994 14530 39006
rect 25342 38994 25394 39006
rect 27582 39058 27634 39070
rect 28702 39058 28754 39070
rect 28354 39006 28366 39058
rect 28418 39006 28430 39058
rect 27582 38994 27634 39006
rect 28702 38994 28754 39006
rect 30382 39058 30434 39070
rect 30382 38994 30434 39006
rect 32510 39058 32562 39070
rect 32510 38994 32562 39006
rect 33966 39058 34018 39070
rect 33966 38994 34018 39006
rect 35646 39058 35698 39070
rect 35646 38994 35698 39006
rect 18622 38946 18674 38958
rect 7298 38894 7310 38946
rect 7362 38894 7374 38946
rect 14690 38894 14702 38946
rect 14754 38894 14766 38946
rect 16706 38894 16718 38946
rect 16770 38894 16782 38946
rect 18622 38882 18674 38894
rect 18846 38946 18898 38958
rect 26910 38946 26962 38958
rect 23874 38894 23886 38946
rect 23938 38894 23950 38946
rect 18846 38882 18898 38894
rect 26910 38882 26962 38894
rect 27022 38946 27074 38958
rect 27022 38882 27074 38894
rect 27246 38946 27298 38958
rect 27246 38882 27298 38894
rect 27470 38946 27522 38958
rect 32062 38946 32114 38958
rect 36094 38946 36146 38958
rect 30930 38894 30942 38946
rect 30994 38894 31006 38946
rect 31490 38894 31502 38946
rect 31554 38894 31566 38946
rect 34514 38894 34526 38946
rect 34578 38894 34590 38946
rect 34962 38894 34974 38946
rect 35026 38894 35038 38946
rect 27470 38882 27522 38894
rect 32062 38882 32114 38894
rect 36094 38882 36146 38894
rect 9886 38834 9938 38846
rect 4274 38782 4286 38834
rect 4338 38782 4350 38834
rect 8082 38782 8094 38834
rect 8146 38782 8158 38834
rect 9886 38770 9938 38782
rect 10558 38834 10610 38846
rect 10558 38770 10610 38782
rect 12126 38834 12178 38846
rect 12126 38770 12178 38782
rect 12462 38834 12514 38846
rect 15262 38834 15314 38846
rect 18510 38834 18562 38846
rect 27694 38834 27746 38846
rect 12786 38782 12798 38834
rect 12850 38782 12862 38834
rect 16034 38782 16046 38834
rect 16098 38782 16110 38834
rect 16482 38782 16494 38834
rect 16546 38782 16558 38834
rect 17490 38782 17502 38834
rect 17554 38782 17566 38834
rect 24658 38782 24670 38834
rect 24722 38782 24734 38834
rect 12462 38770 12514 38782
rect 15262 38770 15314 38782
rect 18510 38770 18562 38782
rect 27694 38770 27746 38782
rect 27918 38834 27970 38846
rect 27918 38770 27970 38782
rect 4846 38722 4898 38734
rect 8542 38722 8594 38734
rect 5170 38670 5182 38722
rect 5234 38670 5246 38722
rect 4846 38658 4898 38670
rect 8542 38658 8594 38670
rect 11454 38722 11506 38734
rect 11454 38658 11506 38670
rect 11902 38722 11954 38734
rect 11902 38658 11954 38670
rect 13582 38722 13634 38734
rect 19182 38722 19234 38734
rect 26574 38722 26626 38734
rect 17826 38670 17838 38722
rect 17890 38670 17902 38722
rect 21746 38670 21758 38722
rect 21810 38670 21822 38722
rect 13582 38658 13634 38670
rect 19182 38658 19234 38670
rect 26574 38658 26626 38670
rect 30718 38722 30770 38734
rect 30718 38658 30770 38670
rect 33294 38722 33346 38734
rect 33294 38658 33346 38670
rect 34302 38722 34354 38734
rect 34302 38658 34354 38670
rect 36654 38722 36706 38734
rect 36654 38658 36706 38670
rect 1934 38610 1986 38622
rect 1934 38546 1986 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 23326 38274 23378 38286
rect 23326 38210 23378 38222
rect 40126 38274 40178 38286
rect 40126 38210 40178 38222
rect 2830 38162 2882 38174
rect 2830 38098 2882 38110
rect 3390 38162 3442 38174
rect 3390 38098 3442 38110
rect 11118 38162 11170 38174
rect 11118 38098 11170 38110
rect 12462 38162 12514 38174
rect 12462 38098 12514 38110
rect 13694 38162 13746 38174
rect 16594 38110 16606 38162
rect 16658 38110 16670 38162
rect 13694 38098 13746 38110
rect 3278 38050 3330 38062
rect 3278 37986 3330 37998
rect 3614 38050 3666 38062
rect 3614 37986 3666 37998
rect 3726 38050 3778 38062
rect 5182 38050 5234 38062
rect 10446 38050 10498 38062
rect 22430 38050 22482 38062
rect 3826 37998 3838 38050
rect 3890 37998 3902 38050
rect 9986 37998 9998 38050
rect 10050 37998 10062 38050
rect 18722 37998 18734 38050
rect 18786 37998 18798 38050
rect 3726 37986 3778 37998
rect 5182 37986 5234 37998
rect 10446 37986 10498 37998
rect 22430 37986 22482 37998
rect 22766 38050 22818 38062
rect 22766 37986 22818 37998
rect 23214 38050 23266 38062
rect 39790 38050 39842 38062
rect 29362 37998 29374 38050
rect 29426 37998 29438 38050
rect 38994 37998 39006 38050
rect 39058 37998 39070 38050
rect 23214 37986 23266 37998
rect 39790 37986 39842 37998
rect 4510 37938 4562 37950
rect 4510 37874 4562 37886
rect 4846 37938 4898 37950
rect 4846 37874 4898 37886
rect 8094 37938 8146 37950
rect 40686 37938 40738 37950
rect 39106 37886 39118 37938
rect 39170 37886 39182 37938
rect 8094 37874 8146 37886
rect 40686 37874 40738 37886
rect 2942 37826 2994 37838
rect 2942 37762 2994 37774
rect 4398 37826 4450 37838
rect 4398 37762 4450 37774
rect 4958 37826 5010 37838
rect 4958 37762 5010 37774
rect 7758 37826 7810 37838
rect 7758 37762 7810 37774
rect 10222 37826 10274 37838
rect 10222 37762 10274 37774
rect 10334 37826 10386 37838
rect 10334 37762 10386 37774
rect 10558 37826 10610 37838
rect 10558 37762 10610 37774
rect 20302 37826 20354 37838
rect 20302 37762 20354 37774
rect 22094 37826 22146 37838
rect 22094 37762 22146 37774
rect 22542 37826 22594 37838
rect 22542 37762 22594 37774
rect 23326 37826 23378 37838
rect 41134 37826 41186 37838
rect 29138 37774 29150 37826
rect 29202 37774 29214 37826
rect 23326 37762 23378 37774
rect 41134 37762 41186 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 7646 37490 7698 37502
rect 7646 37426 7698 37438
rect 9438 37490 9490 37502
rect 9438 37426 9490 37438
rect 11902 37490 11954 37502
rect 11902 37426 11954 37438
rect 13806 37490 13858 37502
rect 13806 37426 13858 37438
rect 18622 37490 18674 37502
rect 28814 37490 28866 37502
rect 19618 37438 19630 37490
rect 19682 37438 19694 37490
rect 18622 37426 18674 37438
rect 28814 37426 28866 37438
rect 29374 37490 29426 37502
rect 29374 37426 29426 37438
rect 32510 37490 32562 37502
rect 32510 37426 32562 37438
rect 34302 37490 34354 37502
rect 34302 37426 34354 37438
rect 34862 37378 34914 37390
rect 9538 37326 9550 37378
rect 9602 37326 9614 37378
rect 11442 37326 11454 37378
rect 11506 37326 11518 37378
rect 12450 37326 12462 37378
rect 12514 37326 12526 37378
rect 14242 37326 14254 37378
rect 14306 37326 14318 37378
rect 16146 37326 16158 37378
rect 16210 37326 16222 37378
rect 17602 37326 17614 37378
rect 17666 37326 17678 37378
rect 18050 37326 18062 37378
rect 18114 37326 18126 37378
rect 27906 37326 27918 37378
rect 27970 37326 27982 37378
rect 28130 37326 28142 37378
rect 28194 37326 28206 37378
rect 33282 37326 33294 37378
rect 33346 37326 33358 37378
rect 33730 37326 33742 37378
rect 33794 37326 33806 37378
rect 34862 37314 34914 37326
rect 5630 37266 5682 37278
rect 2370 37214 2382 37266
rect 2434 37214 2446 37266
rect 5630 37202 5682 37214
rect 7982 37266 8034 37278
rect 28478 37266 28530 37278
rect 9874 37214 9886 37266
rect 9938 37214 9950 37266
rect 10658 37214 10670 37266
rect 10722 37214 10734 37266
rect 10882 37214 10894 37266
rect 10946 37214 10958 37266
rect 12674 37214 12686 37266
rect 12738 37214 12750 37266
rect 14802 37214 14814 37266
rect 14866 37214 14878 37266
rect 15362 37214 15374 37266
rect 15426 37214 15438 37266
rect 15810 37214 15822 37266
rect 15874 37214 15886 37266
rect 7982 37202 8034 37214
rect 28478 37202 28530 37214
rect 29934 37266 29986 37278
rect 29934 37202 29986 37214
rect 13246 37154 13298 37166
rect 16830 37154 16882 37166
rect 3042 37102 3054 37154
rect 3106 37102 3118 37154
rect 5170 37102 5182 37154
rect 5234 37102 5246 37154
rect 14466 37102 14478 37154
rect 14530 37102 14542 37154
rect 13246 37090 13298 37102
rect 16830 37090 16882 37102
rect 19070 37154 19122 37166
rect 19070 37090 19122 37102
rect 20078 37154 20130 37166
rect 20078 37090 20130 37102
rect 20526 37154 20578 37166
rect 20526 37090 20578 37102
rect 27246 37154 27298 37166
rect 27246 37090 27298 37102
rect 33966 37154 34018 37166
rect 33966 37090 34018 37102
rect 35422 37154 35474 37166
rect 35422 37090 35474 37102
rect 18286 37042 18338 37054
rect 18286 36978 18338 36990
rect 19294 37042 19346 37054
rect 19294 36978 19346 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 4958 36706 5010 36718
rect 4958 36642 5010 36654
rect 12014 36706 12066 36718
rect 12014 36642 12066 36654
rect 1934 36594 1986 36606
rect 1934 36530 1986 36542
rect 5742 36594 5794 36606
rect 12238 36594 12290 36606
rect 15598 36594 15650 36606
rect 20302 36594 20354 36606
rect 11106 36542 11118 36594
rect 11170 36542 11182 36594
rect 13570 36542 13582 36594
rect 13634 36542 13646 36594
rect 19282 36542 19294 36594
rect 19346 36542 19358 36594
rect 5742 36530 5794 36542
rect 12238 36530 12290 36542
rect 15598 36530 15650 36542
rect 20302 36530 20354 36542
rect 20862 36594 20914 36606
rect 20862 36530 20914 36542
rect 21422 36594 21474 36606
rect 32610 36542 32622 36594
rect 32674 36542 32686 36594
rect 21422 36530 21474 36542
rect 5630 36482 5682 36494
rect 6078 36482 6130 36494
rect 8878 36482 8930 36494
rect 9774 36482 9826 36494
rect 4274 36430 4286 36482
rect 4338 36430 4350 36482
rect 5842 36430 5854 36482
rect 5906 36430 5918 36482
rect 6402 36430 6414 36482
rect 6466 36430 6478 36482
rect 9538 36430 9550 36482
rect 9602 36430 9614 36482
rect 5630 36418 5682 36430
rect 6078 36418 6130 36430
rect 8878 36418 8930 36430
rect 9774 36418 9826 36430
rect 9998 36482 10050 36494
rect 12462 36482 12514 36494
rect 13694 36482 13746 36494
rect 11554 36430 11566 36482
rect 11618 36430 11630 36482
rect 13458 36430 13470 36482
rect 13522 36430 13534 36482
rect 9998 36418 10050 36430
rect 12462 36418 12514 36430
rect 13694 36418 13746 36430
rect 13918 36482 13970 36494
rect 13918 36418 13970 36430
rect 14030 36482 14082 36494
rect 18398 36482 18450 36494
rect 15138 36430 15150 36482
rect 15202 36430 15214 36482
rect 16594 36430 16606 36482
rect 16658 36430 16670 36482
rect 17154 36430 17166 36482
rect 17218 36430 17230 36482
rect 17378 36430 17390 36482
rect 17442 36430 17454 36482
rect 30034 36430 30046 36482
rect 30098 36430 30110 36482
rect 41010 36430 41022 36482
rect 41074 36430 41086 36482
rect 14030 36418 14082 36430
rect 18398 36418 18450 36430
rect 5070 36370 5122 36382
rect 5070 36306 5122 36318
rect 8206 36370 8258 36382
rect 8206 36306 8258 36318
rect 8430 36370 8482 36382
rect 8430 36306 8482 36318
rect 10222 36370 10274 36382
rect 22206 36370 22258 36382
rect 11778 36318 11790 36370
rect 11842 36318 11854 36370
rect 16146 36318 16158 36370
rect 16210 36318 16222 36370
rect 17938 36318 17950 36370
rect 18002 36318 18014 36370
rect 10222 36306 10274 36318
rect 22206 36306 22258 36318
rect 22318 36370 22370 36382
rect 22318 36306 22370 36318
rect 47630 36370 47682 36382
rect 47630 36306 47682 36318
rect 48190 36370 48242 36382
rect 48190 36306 48242 36318
rect 6862 36258 6914 36270
rect 6862 36194 6914 36206
rect 8654 36258 8706 36270
rect 8654 36194 8706 36206
rect 9886 36258 9938 36270
rect 9886 36194 9938 36206
rect 10670 36258 10722 36270
rect 10670 36194 10722 36206
rect 12014 36258 12066 36270
rect 12014 36194 12066 36206
rect 12910 36258 12962 36270
rect 12910 36194 12962 36206
rect 14702 36258 14754 36270
rect 14702 36194 14754 36206
rect 15934 36258 15986 36270
rect 15934 36194 15986 36206
rect 18846 36258 18898 36270
rect 18846 36194 18898 36206
rect 19854 36258 19906 36270
rect 19854 36194 19906 36206
rect 21534 36258 21586 36270
rect 21534 36194 21586 36206
rect 22542 36258 22594 36270
rect 22542 36194 22594 36206
rect 22878 36258 22930 36270
rect 22878 36194 22930 36206
rect 28590 36258 28642 36270
rect 47854 36258 47906 36270
rect 41234 36206 41246 36258
rect 41298 36206 41310 36258
rect 28590 36194 28642 36206
rect 47854 36194 47906 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 14814 35922 14866 35934
rect 4610 35870 4622 35922
rect 4674 35870 4686 35922
rect 9538 35870 9550 35922
rect 9602 35870 9614 35922
rect 14814 35858 14866 35870
rect 15710 35922 15762 35934
rect 15710 35858 15762 35870
rect 16046 35922 16098 35934
rect 19182 35922 19234 35934
rect 16370 35870 16382 35922
rect 16434 35870 16446 35922
rect 16046 35858 16098 35870
rect 19182 35858 19234 35870
rect 24558 35922 24610 35934
rect 24558 35858 24610 35870
rect 19294 35810 19346 35822
rect 18610 35758 18622 35810
rect 18674 35758 18686 35810
rect 19294 35746 19346 35758
rect 19742 35810 19794 35822
rect 19742 35746 19794 35758
rect 32174 35810 32226 35822
rect 32174 35746 32226 35758
rect 32398 35810 32450 35822
rect 32398 35746 32450 35758
rect 4958 35698 5010 35710
rect 4274 35646 4286 35698
rect 4338 35646 4350 35698
rect 4958 35634 5010 35646
rect 9886 35698 9938 35710
rect 9886 35634 9938 35646
rect 12350 35698 12402 35710
rect 12350 35634 12402 35646
rect 14030 35698 14082 35710
rect 14030 35634 14082 35646
rect 14366 35698 14418 35710
rect 14366 35634 14418 35646
rect 18286 35698 18338 35710
rect 24098 35646 24110 35698
rect 24162 35646 24174 35698
rect 33058 35646 33070 35698
rect 33122 35646 33134 35698
rect 36418 35646 36430 35698
rect 36482 35646 36494 35698
rect 18286 35634 18338 35646
rect 10446 35586 10498 35598
rect 10446 35522 10498 35534
rect 12574 35586 12626 35598
rect 12574 35522 12626 35534
rect 15262 35586 15314 35598
rect 15262 35522 15314 35534
rect 17502 35586 17554 35598
rect 17502 35522 17554 35534
rect 18062 35586 18114 35598
rect 18062 35522 18114 35534
rect 18846 35586 18898 35598
rect 18846 35522 18898 35534
rect 19070 35586 19122 35598
rect 29822 35586 29874 35598
rect 21186 35534 21198 35586
rect 21250 35534 21262 35586
rect 23314 35534 23326 35586
rect 23378 35534 23390 35586
rect 19070 35522 19122 35534
rect 29822 35522 29874 35534
rect 31838 35586 31890 35598
rect 32498 35534 32510 35586
rect 32562 35534 32574 35586
rect 33842 35534 33854 35586
rect 33906 35534 33918 35586
rect 35970 35534 35982 35586
rect 36034 35534 36046 35586
rect 37202 35534 37214 35586
rect 37266 35534 37278 35586
rect 39330 35534 39342 35586
rect 39394 35534 39406 35586
rect 31838 35522 31890 35534
rect 1934 35474 1986 35486
rect 12002 35422 12014 35474
rect 12066 35422 12078 35474
rect 1934 35410 1986 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 4734 35138 4786 35150
rect 4734 35074 4786 35086
rect 7310 35138 7362 35150
rect 34750 35138 34802 35150
rect 24882 35086 24894 35138
rect 24946 35086 24958 35138
rect 30594 35086 30606 35138
rect 30658 35086 30670 35138
rect 7310 35074 7362 35086
rect 34750 35074 34802 35086
rect 41246 35138 41298 35150
rect 41246 35074 41298 35086
rect 41582 35138 41634 35150
rect 41582 35074 41634 35086
rect 8318 35026 8370 35038
rect 30270 35026 30322 35038
rect 13682 34974 13694 35026
rect 13746 34974 13758 35026
rect 8318 34962 8370 34974
rect 30270 34962 30322 34974
rect 32734 35026 32786 35038
rect 32734 34962 32786 34974
rect 36094 35026 36146 35038
rect 36094 34962 36146 34974
rect 2830 34914 2882 34926
rect 3614 34914 3666 34926
rect 4062 34914 4114 34926
rect 3266 34862 3278 34914
rect 3330 34862 3342 34914
rect 3826 34862 3838 34914
rect 3890 34862 3902 34914
rect 2830 34850 2882 34862
rect 3614 34850 3666 34862
rect 4062 34850 4114 34862
rect 8990 34914 9042 34926
rect 8990 34850 9042 34862
rect 9774 34914 9826 34926
rect 22430 34914 22482 34926
rect 24334 34914 24386 34926
rect 12226 34862 12238 34914
rect 12290 34862 12302 34914
rect 18722 34862 18734 34914
rect 18786 34862 18798 34914
rect 22866 34862 22878 34914
rect 22930 34862 22942 34914
rect 9774 34850 9826 34862
rect 22430 34850 22482 34862
rect 24334 34850 24386 34862
rect 24558 34914 24610 34926
rect 24558 34850 24610 34862
rect 30046 34914 30098 34926
rect 35074 34862 35086 34914
rect 35138 34862 35150 34914
rect 40450 34862 40462 34914
rect 40514 34862 40526 34914
rect 30046 34850 30098 34862
rect 2942 34802 2994 34814
rect 2942 34738 2994 34750
rect 4398 34802 4450 34814
rect 4398 34738 4450 34750
rect 5630 34802 5682 34814
rect 5630 34738 5682 34750
rect 5966 34802 6018 34814
rect 5966 34738 6018 34750
rect 7310 34802 7362 34814
rect 7310 34738 7362 34750
rect 7422 34802 7474 34814
rect 7422 34738 7474 34750
rect 9438 34802 9490 34814
rect 12574 34802 12626 34814
rect 9650 34750 9662 34802
rect 9714 34750 9726 34802
rect 9438 34738 9490 34750
rect 12574 34738 12626 34750
rect 29150 34802 29202 34814
rect 29150 34738 29202 34750
rect 29710 34802 29762 34814
rect 42142 34802 42194 34814
rect 40674 34750 40686 34802
rect 40738 34750 40750 34802
rect 29710 34738 29762 34750
rect 42142 34738 42194 34750
rect 2382 34690 2434 34702
rect 2382 34626 2434 34638
rect 2718 34690 2770 34702
rect 4622 34690 4674 34702
rect 3602 34638 3614 34690
rect 3666 34638 3678 34690
rect 2718 34626 2770 34638
rect 4622 34626 4674 34638
rect 7870 34690 7922 34702
rect 7870 34626 7922 34638
rect 8766 34690 8818 34702
rect 8766 34626 8818 34638
rect 12462 34690 12514 34702
rect 12462 34626 12514 34638
rect 12686 34690 12738 34702
rect 12686 34626 12738 34638
rect 12798 34690 12850 34702
rect 12798 34626 12850 34638
rect 19182 34690 19234 34702
rect 19182 34626 19234 34638
rect 22878 34690 22930 34702
rect 22878 34626 22930 34638
rect 29262 34690 29314 34702
rect 29262 34626 29314 34638
rect 34862 34690 34914 34702
rect 34862 34626 34914 34638
rect 40126 34690 40178 34702
rect 40126 34626 40178 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 2046 34354 2098 34366
rect 2046 34290 2098 34302
rect 13134 34354 13186 34366
rect 18510 34354 18562 34366
rect 13458 34302 13470 34354
rect 13522 34302 13534 34354
rect 13134 34290 13186 34302
rect 18510 34290 18562 34302
rect 25342 34354 25394 34366
rect 25342 34290 25394 34302
rect 35534 34354 35586 34366
rect 35534 34290 35586 34302
rect 3838 34242 3890 34254
rect 3838 34178 3890 34190
rect 4062 34242 4114 34254
rect 4062 34178 4114 34190
rect 12238 34242 12290 34254
rect 12238 34178 12290 34190
rect 12350 34242 12402 34254
rect 12350 34178 12402 34190
rect 14030 34242 14082 34254
rect 19518 34242 19570 34254
rect 19282 34190 19294 34242
rect 19346 34190 19358 34242
rect 14030 34178 14082 34190
rect 19518 34178 19570 34190
rect 26126 34242 26178 34254
rect 26126 34178 26178 34190
rect 26462 34242 26514 34254
rect 26462 34178 26514 34190
rect 1710 34130 1762 34142
rect 12462 34130 12514 34142
rect 12002 34078 12014 34130
rect 12066 34078 12078 34130
rect 1710 34066 1762 34078
rect 12462 34066 12514 34078
rect 13918 34130 13970 34142
rect 18622 34130 18674 34142
rect 14242 34078 14254 34130
rect 14306 34078 14318 34130
rect 13918 34066 13970 34078
rect 18622 34066 18674 34078
rect 19070 34130 19122 34142
rect 35198 34130 35250 34142
rect 24434 34078 24446 34130
rect 24498 34078 24510 34130
rect 30370 34078 30382 34130
rect 30434 34078 30446 34130
rect 19070 34066 19122 34078
rect 35198 34066 35250 34078
rect 35534 34130 35586 34142
rect 35534 34066 35586 34078
rect 35870 34130 35922 34142
rect 35870 34066 35922 34078
rect 2494 34018 2546 34030
rect 2494 33954 2546 33966
rect 3390 34018 3442 34030
rect 4510 34018 4562 34030
rect 3714 33966 3726 34018
rect 3778 33966 3790 34018
rect 3390 33954 3442 33966
rect 4510 33954 4562 33966
rect 4958 34018 5010 34030
rect 4958 33954 5010 33966
rect 18846 34018 18898 34030
rect 18846 33954 18898 33966
rect 19966 34018 20018 34030
rect 30942 34018 30994 34030
rect 21634 33966 21646 34018
rect 21698 33966 21710 34018
rect 23762 33966 23774 34018
rect 23826 33966 23838 34018
rect 26898 33966 26910 34018
rect 26962 33966 26974 34018
rect 27458 33966 27470 34018
rect 27522 33966 27534 34018
rect 29586 33966 29598 34018
rect 29650 33966 29662 34018
rect 19966 33954 20018 33966
rect 30942 33954 30994 33966
rect 11566 33906 11618 33918
rect 4274 33854 4286 33906
rect 4338 33903 4350 33906
rect 4610 33903 4622 33906
rect 4338 33857 4622 33903
rect 4338 33854 4350 33857
rect 4610 33854 4622 33857
rect 4674 33903 4686 33906
rect 4946 33903 4958 33906
rect 4674 33857 4958 33903
rect 4674 33854 4686 33857
rect 4946 33854 4958 33857
rect 5010 33854 5022 33906
rect 30594 33854 30606 33906
rect 30658 33903 30670 33906
rect 30930 33903 30942 33906
rect 30658 33857 30942 33903
rect 30658 33854 30670 33857
rect 30930 33854 30942 33857
rect 30994 33854 31006 33906
rect 11566 33842 11618 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 23102 33570 23154 33582
rect 34974 33570 35026 33582
rect 34178 33518 34190 33570
rect 34242 33567 34254 33570
rect 34514 33567 34526 33570
rect 34242 33521 34526 33567
rect 34242 33518 34254 33521
rect 34514 33518 34526 33521
rect 34578 33518 34590 33570
rect 23102 33506 23154 33518
rect 34974 33506 35026 33518
rect 17726 33458 17778 33470
rect 17726 33394 17778 33406
rect 27022 33458 27074 33470
rect 27022 33394 27074 33406
rect 28590 33458 28642 33470
rect 28590 33394 28642 33406
rect 29262 33458 29314 33470
rect 29262 33394 29314 33406
rect 34526 33458 34578 33470
rect 34526 33394 34578 33406
rect 35534 33458 35586 33470
rect 38882 33406 38894 33458
rect 38946 33406 38958 33458
rect 41010 33406 41022 33458
rect 41074 33406 41086 33458
rect 35534 33394 35586 33406
rect 9550 33346 9602 33358
rect 9550 33282 9602 33294
rect 17838 33346 17890 33358
rect 17838 33282 17890 33294
rect 18510 33346 18562 33358
rect 18510 33282 18562 33294
rect 27694 33346 27746 33358
rect 27694 33282 27746 33294
rect 29038 33346 29090 33358
rect 29038 33282 29090 33294
rect 29374 33346 29426 33358
rect 35310 33346 35362 33358
rect 30146 33294 30158 33346
rect 30210 33294 30222 33346
rect 29374 33282 29426 33294
rect 35310 33282 35362 33294
rect 35870 33346 35922 33358
rect 38098 33294 38110 33346
rect 38162 33294 38174 33346
rect 35870 33282 35922 33294
rect 9774 33234 9826 33246
rect 9774 33170 9826 33182
rect 9886 33234 9938 33246
rect 9886 33170 9938 33182
rect 17054 33234 17106 33246
rect 17054 33170 17106 33182
rect 17390 33234 17442 33246
rect 17390 33170 17442 33182
rect 22990 33234 23042 33246
rect 22990 33170 23042 33182
rect 27358 33234 27410 33246
rect 27358 33170 27410 33182
rect 27470 33234 27522 33246
rect 27470 33170 27522 33182
rect 27918 33234 27970 33246
rect 27918 33170 27970 33182
rect 28030 33234 28082 33246
rect 28030 33170 28082 33182
rect 28254 33234 28306 33246
rect 28254 33170 28306 33182
rect 29710 33234 29762 33246
rect 29710 33170 29762 33182
rect 30382 33234 30434 33246
rect 35758 33234 35810 33246
rect 30382 33170 30434 33182
rect 34862 33178 34914 33190
rect 10446 33122 10498 33134
rect 10446 33058 10498 33070
rect 12910 33122 12962 33134
rect 12910 33058 12962 33070
rect 17614 33122 17666 33134
rect 17614 33058 17666 33070
rect 17950 33122 18002 33134
rect 17950 33058 18002 33070
rect 22654 33122 22706 33134
rect 35758 33170 35810 33182
rect 34862 33114 34914 33126
rect 34974 33122 35026 33134
rect 22654 33058 22706 33070
rect 34974 33058 35026 33070
rect 37774 33122 37826 33134
rect 37774 33058 37826 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 19518 32786 19570 32798
rect 12002 32734 12014 32786
rect 12066 32734 12078 32786
rect 13234 32734 13246 32786
rect 13298 32734 13310 32786
rect 19518 32722 19570 32734
rect 26574 32786 26626 32798
rect 26574 32722 26626 32734
rect 28366 32786 28418 32798
rect 28366 32722 28418 32734
rect 29374 32786 29426 32798
rect 29374 32722 29426 32734
rect 35086 32786 35138 32798
rect 35086 32722 35138 32734
rect 10670 32674 10722 32686
rect 10670 32610 10722 32622
rect 18174 32674 18226 32686
rect 18174 32610 18226 32622
rect 18286 32674 18338 32686
rect 18286 32610 18338 32622
rect 27022 32674 27074 32686
rect 27022 32610 27074 32622
rect 27470 32674 27522 32686
rect 27470 32610 27522 32622
rect 27582 32674 27634 32686
rect 27582 32610 27634 32622
rect 29150 32674 29202 32686
rect 29150 32610 29202 32622
rect 34862 32674 34914 32686
rect 34862 32610 34914 32622
rect 35422 32674 35474 32686
rect 35422 32610 35474 32622
rect 35646 32674 35698 32686
rect 35646 32610 35698 32622
rect 11006 32562 11058 32574
rect 4274 32510 4286 32562
rect 4338 32510 4350 32562
rect 11006 32498 11058 32510
rect 12350 32562 12402 32574
rect 12350 32498 12402 32510
rect 12910 32562 12962 32574
rect 12910 32498 12962 32510
rect 13806 32562 13858 32574
rect 13806 32498 13858 32510
rect 14366 32562 14418 32574
rect 14366 32498 14418 32510
rect 18062 32562 18114 32574
rect 18062 32498 18114 32510
rect 27134 32562 27186 32574
rect 27134 32498 27186 32510
rect 27806 32562 27858 32574
rect 27806 32498 27858 32510
rect 28030 32562 28082 32574
rect 28030 32498 28082 32510
rect 28366 32562 28418 32574
rect 28366 32498 28418 32510
rect 28702 32562 28754 32574
rect 28702 32498 28754 32510
rect 29038 32562 29090 32574
rect 29038 32498 29090 32510
rect 34750 32562 34802 32574
rect 34750 32498 34802 32510
rect 35310 32562 35362 32574
rect 35310 32498 35362 32510
rect 35870 32562 35922 32574
rect 35870 32498 35922 32510
rect 36094 32562 36146 32574
rect 36094 32498 36146 32510
rect 36430 32562 36482 32574
rect 37426 32510 37438 32562
rect 37490 32510 37502 32562
rect 36430 32498 36482 32510
rect 5070 32450 5122 32462
rect 5070 32386 5122 32398
rect 12574 32450 12626 32462
rect 12574 32386 12626 32398
rect 20302 32450 20354 32462
rect 20302 32386 20354 32398
rect 29710 32450 29762 32462
rect 29710 32386 29762 32398
rect 34414 32450 34466 32462
rect 34414 32386 34466 32398
rect 36318 32450 36370 32462
rect 36318 32386 36370 32398
rect 36878 32450 36930 32462
rect 38210 32398 38222 32450
rect 38274 32398 38286 32450
rect 40338 32398 40350 32450
rect 40402 32398 40414 32450
rect 36878 32386 36930 32398
rect 1934 32338 1986 32350
rect 27022 32338 27074 32350
rect 17602 32286 17614 32338
rect 17666 32286 17678 32338
rect 29474 32286 29486 32338
rect 29538 32335 29550 32338
rect 29810 32335 29822 32338
rect 29538 32289 29822 32335
rect 29538 32286 29550 32289
rect 29810 32286 29822 32289
rect 29874 32286 29886 32338
rect 1934 32274 1986 32286
rect 27022 32274 27074 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 12574 32002 12626 32014
rect 12574 31938 12626 31950
rect 9102 31890 9154 31902
rect 1922 31838 1934 31890
rect 1986 31838 1998 31890
rect 9102 31826 9154 31838
rect 9886 31890 9938 31902
rect 9886 31826 9938 31838
rect 10110 31890 10162 31902
rect 10110 31826 10162 31838
rect 10782 31890 10834 31902
rect 10782 31826 10834 31838
rect 14926 31890 14978 31902
rect 30830 31890 30882 31902
rect 19394 31838 19406 31890
rect 19458 31838 19470 31890
rect 14926 31826 14978 31838
rect 30830 31826 30882 31838
rect 5742 31778 5794 31790
rect 4834 31726 4846 31778
rect 4898 31726 4910 31778
rect 5742 31714 5794 31726
rect 8878 31778 8930 31790
rect 8878 31714 8930 31726
rect 9326 31778 9378 31790
rect 9326 31714 9378 31726
rect 10334 31778 10386 31790
rect 10334 31714 10386 31726
rect 12126 31778 12178 31790
rect 12126 31714 12178 31726
rect 19742 31778 19794 31790
rect 19954 31726 19966 31778
rect 20018 31726 20030 31778
rect 31154 31726 31166 31778
rect 31218 31726 31230 31778
rect 19742 31714 19794 31726
rect 11902 31666 11954 31678
rect 4050 31614 4062 31666
rect 4114 31614 4126 31666
rect 9650 31614 9662 31666
rect 9714 31614 9726 31666
rect 11902 31602 11954 31614
rect 12014 31666 12066 31678
rect 12014 31602 12066 31614
rect 12686 31666 12738 31678
rect 27234 31614 27246 31666
rect 27298 31614 27310 31666
rect 34402 31614 34414 31666
rect 34466 31614 34478 31666
rect 12686 31602 12738 31614
rect 5854 31554 5906 31566
rect 5854 31490 5906 31502
rect 8318 31554 8370 31566
rect 13582 31554 13634 31566
rect 8530 31502 8542 31554
rect 8594 31502 8606 31554
rect 9762 31502 9774 31554
rect 9826 31502 9838 31554
rect 11442 31502 11454 31554
rect 11506 31502 11518 31554
rect 8318 31490 8370 31502
rect 13582 31490 13634 31502
rect 19070 31554 19122 31566
rect 19070 31490 19122 31502
rect 19406 31554 19458 31566
rect 19406 31490 19458 31502
rect 19518 31554 19570 31566
rect 19518 31490 19570 31502
rect 20526 31554 20578 31566
rect 20526 31490 20578 31502
rect 27582 31554 27634 31566
rect 27582 31490 27634 31502
rect 37102 31554 37154 31566
rect 37102 31490 37154 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 7982 31218 8034 31230
rect 7982 31154 8034 31166
rect 9438 31218 9490 31230
rect 9438 31154 9490 31166
rect 10894 31218 10946 31230
rect 10894 31154 10946 31166
rect 14590 31218 14642 31230
rect 14590 31154 14642 31166
rect 18958 31218 19010 31230
rect 18958 31154 19010 31166
rect 19070 31218 19122 31230
rect 19070 31154 19122 31166
rect 19182 31218 19234 31230
rect 19182 31154 19234 31166
rect 19966 31218 20018 31230
rect 19966 31154 20018 31166
rect 22766 31218 22818 31230
rect 22766 31154 22818 31166
rect 23214 31218 23266 31230
rect 23214 31154 23266 31166
rect 24446 31218 24498 31230
rect 24446 31154 24498 31166
rect 28030 31218 28082 31230
rect 28030 31154 28082 31166
rect 33742 31218 33794 31230
rect 33742 31154 33794 31166
rect 34190 31218 34242 31230
rect 34190 31154 34242 31166
rect 35870 31218 35922 31230
rect 35870 31154 35922 31166
rect 36206 31218 36258 31230
rect 36206 31154 36258 31166
rect 36990 31218 37042 31230
rect 36990 31154 37042 31166
rect 37998 31218 38050 31230
rect 37998 31154 38050 31166
rect 41246 31218 41298 31230
rect 41246 31154 41298 31166
rect 41694 31218 41746 31230
rect 41694 31154 41746 31166
rect 43486 31218 43538 31230
rect 43486 31154 43538 31166
rect 8094 31106 8146 31118
rect 14478 31106 14530 31118
rect 6066 31054 6078 31106
rect 6130 31054 6142 31106
rect 13794 31054 13806 31106
rect 13858 31054 13870 31106
rect 8094 31042 8146 31054
rect 14478 31042 14530 31054
rect 15262 31106 15314 31118
rect 15262 31042 15314 31054
rect 15374 31106 15426 31118
rect 27246 31106 27298 31118
rect 18162 31054 18174 31106
rect 18226 31054 18238 31106
rect 20290 31054 20302 31106
rect 20354 31054 20366 31106
rect 22306 31054 22318 31106
rect 22370 31054 22382 31106
rect 15374 31042 15426 31054
rect 27246 31042 27298 31054
rect 27358 31106 27410 31118
rect 27358 31042 27410 31054
rect 27582 31106 27634 31118
rect 27582 31042 27634 31054
rect 28366 31106 28418 31118
rect 28366 31042 28418 31054
rect 28814 31106 28866 31118
rect 28814 31042 28866 31054
rect 28926 31106 28978 31118
rect 28926 31042 28978 31054
rect 34078 31106 34130 31118
rect 36430 31106 36482 31118
rect 34850 31054 34862 31106
rect 34914 31054 34926 31106
rect 34078 31042 34130 31054
rect 36430 31042 36482 31054
rect 36878 31106 36930 31118
rect 47854 31106 47906 31118
rect 42578 31054 42590 31106
rect 42642 31054 42654 31106
rect 36878 31042 36930 31054
rect 47854 31042 47906 31054
rect 7310 30994 7362 31006
rect 6738 30942 6750 30994
rect 6802 30942 6814 30994
rect 7310 30930 7362 30942
rect 7758 30994 7810 31006
rect 9102 30994 9154 31006
rect 8754 30942 8766 30994
rect 8818 30942 8830 30994
rect 7758 30930 7810 30942
rect 9102 30930 9154 30942
rect 9550 30994 9602 31006
rect 9550 30930 9602 30942
rect 9774 30994 9826 31006
rect 9774 30930 9826 30942
rect 9998 30994 10050 31006
rect 10558 30994 10610 31006
rect 14030 30994 14082 31006
rect 19294 30994 19346 31006
rect 20750 30994 20802 31006
rect 27694 30994 27746 31006
rect 10210 30942 10222 30994
rect 10274 30942 10286 30994
rect 13570 30942 13582 30994
rect 13634 30942 13646 30994
rect 15586 30942 15598 30994
rect 15650 30942 15662 30994
rect 18386 30942 18398 30994
rect 18450 30942 18462 30994
rect 19506 30942 19518 30994
rect 19570 30942 19582 30994
rect 20626 30942 20638 30994
rect 20690 30942 20702 30994
rect 21522 30942 21534 30994
rect 21586 30942 21598 30994
rect 21746 30942 21758 30994
rect 21810 30942 21822 30994
rect 9998 30930 10050 30942
rect 10558 30930 10610 30942
rect 14030 30930 14082 30942
rect 19294 30930 19346 30942
rect 20750 30930 20802 30942
rect 27694 30930 27746 30942
rect 28142 30994 28194 31006
rect 28142 30930 28194 30942
rect 28590 30994 28642 31006
rect 36542 30994 36594 31006
rect 43150 30994 43202 31006
rect 34738 30942 34750 30994
rect 34802 30942 34814 30994
rect 42354 30942 42366 30994
rect 42418 30942 42430 30994
rect 28590 30930 28642 30942
rect 36542 30930 36594 30942
rect 43150 30930 43202 30942
rect 48190 30994 48242 31006
rect 48190 30930 48242 30942
rect 7646 30882 7698 30894
rect 3938 30830 3950 30882
rect 4002 30830 4014 30882
rect 7646 30818 7698 30830
rect 8318 30882 8370 30894
rect 8318 30818 8370 30830
rect 8542 30882 8594 30894
rect 8542 30818 8594 30830
rect 11454 30882 11506 30894
rect 11454 30818 11506 30830
rect 13246 30882 13298 30894
rect 13246 30818 13298 30830
rect 14254 30882 14306 30894
rect 14254 30818 14306 30830
rect 16046 30882 16098 30894
rect 16046 30818 16098 30830
rect 17838 30882 17890 30894
rect 17838 30818 17890 30830
rect 29374 30882 29426 30894
rect 29374 30818 29426 30830
rect 37550 30882 37602 30894
rect 37550 30818 37602 30830
rect 47630 30882 47682 30894
rect 47630 30818 47682 30830
rect 34190 30770 34242 30782
rect 10658 30718 10670 30770
rect 10722 30767 10734 30770
rect 11442 30767 11454 30770
rect 10722 30721 11454 30767
rect 10722 30718 10734 30721
rect 11442 30718 11454 30721
rect 11506 30718 11518 30770
rect 14802 30718 14814 30770
rect 14866 30718 14878 30770
rect 34190 30706 34242 30718
rect 35534 30770 35586 30782
rect 35534 30706 35586 30718
rect 36990 30770 37042 30782
rect 36990 30706 37042 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 25230 30434 25282 30446
rect 25230 30370 25282 30382
rect 1934 30322 1986 30334
rect 1934 30258 1986 30270
rect 18510 30322 18562 30334
rect 18510 30258 18562 30270
rect 19742 30322 19794 30334
rect 19742 30258 19794 30270
rect 20638 30322 20690 30334
rect 34414 30322 34466 30334
rect 21634 30270 21646 30322
rect 21698 30270 21710 30322
rect 33954 30270 33966 30322
rect 34018 30270 34030 30322
rect 41794 30270 41806 30322
rect 41858 30270 41870 30322
rect 20638 30258 20690 30270
rect 34414 30258 34466 30270
rect 9102 30210 9154 30222
rect 3938 30158 3950 30210
rect 4002 30158 4014 30210
rect 9102 30146 9154 30158
rect 9774 30210 9826 30222
rect 9774 30146 9826 30158
rect 14254 30210 14306 30222
rect 25006 30210 25058 30222
rect 26014 30210 26066 30222
rect 14690 30158 14702 30210
rect 14754 30158 14766 30210
rect 15586 30158 15598 30210
rect 15650 30158 15662 30210
rect 16706 30158 16718 30210
rect 16770 30158 16782 30210
rect 24546 30158 24558 30210
rect 24610 30158 24622 30210
rect 25554 30158 25566 30210
rect 25618 30158 25630 30210
rect 14254 30146 14306 30158
rect 25006 30146 25058 30158
rect 26014 30146 26066 30158
rect 30158 30210 30210 30222
rect 30158 30146 30210 30158
rect 30382 30210 30434 30222
rect 35982 30210 36034 30222
rect 31154 30158 31166 30210
rect 31218 30158 31230 30210
rect 31826 30158 31838 30210
rect 31890 30158 31902 30210
rect 38882 30158 38894 30210
rect 38946 30158 38958 30210
rect 30382 30146 30434 30158
rect 35982 30146 36034 30158
rect 10222 30098 10274 30110
rect 35310 30098 35362 30110
rect 8754 30046 8766 30098
rect 8818 30046 8830 30098
rect 9426 30046 9438 30098
rect 9490 30046 9502 30098
rect 15698 30046 15710 30098
rect 15762 30046 15774 30098
rect 16594 30046 16606 30098
rect 16658 30046 16670 30098
rect 23762 30046 23774 30098
rect 23826 30046 23838 30098
rect 30706 30046 30718 30098
rect 30770 30046 30782 30098
rect 10222 30034 10274 30046
rect 35310 30034 35362 30046
rect 35534 30098 35586 30110
rect 35534 30034 35586 30046
rect 35758 30098 35810 30110
rect 39666 30046 39678 30098
rect 39730 30046 39742 30098
rect 35758 30034 35810 30046
rect 14478 29986 14530 29998
rect 14478 29922 14530 29934
rect 17614 29986 17666 29998
rect 17614 29922 17666 29934
rect 17950 29986 18002 29998
rect 17950 29922 18002 29934
rect 19182 29986 19234 29998
rect 19182 29922 19234 29934
rect 20078 29986 20130 29998
rect 20078 29922 20130 29934
rect 35086 29986 35138 29998
rect 35086 29922 35138 29934
rect 36318 29986 36370 29998
rect 36318 29922 36370 29934
rect 38558 29986 38610 29998
rect 38558 29922 38610 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 16046 29650 16098 29662
rect 16046 29586 16098 29598
rect 16718 29650 16770 29662
rect 16718 29586 16770 29598
rect 18510 29650 18562 29662
rect 18510 29586 18562 29598
rect 19406 29650 19458 29662
rect 19406 29586 19458 29598
rect 30942 29650 30994 29662
rect 35198 29650 35250 29662
rect 33506 29598 33518 29650
rect 33570 29598 33582 29650
rect 30942 29586 30994 29598
rect 35198 29586 35250 29598
rect 13694 29538 13746 29550
rect 15934 29538 15986 29550
rect 15138 29486 15150 29538
rect 15202 29486 15214 29538
rect 13694 29474 13746 29486
rect 15934 29474 15986 29486
rect 19966 29538 20018 29550
rect 34862 29538 34914 29550
rect 28354 29486 28366 29538
rect 28418 29486 28430 29538
rect 19966 29474 20018 29486
rect 34862 29474 34914 29486
rect 34974 29538 35026 29550
rect 34974 29474 35026 29486
rect 16270 29426 16322 29438
rect 4274 29374 4286 29426
rect 4338 29374 4350 29426
rect 14018 29374 14030 29426
rect 14082 29374 14094 29426
rect 14802 29374 14814 29426
rect 14866 29374 14878 29426
rect 16270 29362 16322 29374
rect 19518 29426 19570 29438
rect 19518 29362 19570 29374
rect 19630 29426 19682 29438
rect 19630 29362 19682 29374
rect 19742 29426 19794 29438
rect 33182 29426 33234 29438
rect 27682 29374 27694 29426
rect 27746 29374 27758 29426
rect 19742 29362 19794 29374
rect 33182 29362 33234 29374
rect 17614 29314 17666 29326
rect 14690 29262 14702 29314
rect 14754 29262 14766 29314
rect 17614 29250 17666 29262
rect 18062 29314 18114 29326
rect 18062 29250 18114 29262
rect 18958 29314 19010 29326
rect 18958 29250 19010 29262
rect 20414 29314 20466 29326
rect 20414 29250 20466 29262
rect 24670 29314 24722 29326
rect 34526 29314 34578 29326
rect 30482 29262 30494 29314
rect 30546 29262 30558 29314
rect 24670 29250 24722 29262
rect 34526 29250 34578 29262
rect 1934 29202 1986 29214
rect 1934 29138 1986 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 14802 28814 14814 28866
rect 14866 28863 14878 28866
rect 15474 28863 15486 28866
rect 14866 28817 15486 28863
rect 14866 28814 14878 28817
rect 15474 28814 15486 28817
rect 15538 28814 15550 28866
rect 5742 28754 5794 28766
rect 2146 28702 2158 28754
rect 2210 28702 2222 28754
rect 5742 28690 5794 28702
rect 7534 28754 7586 28766
rect 7534 28690 7586 28702
rect 8990 28754 9042 28766
rect 35982 28754 36034 28766
rect 35074 28702 35086 28754
rect 35138 28702 35150 28754
rect 8990 28690 9042 28702
rect 35982 28690 36034 28702
rect 39566 28754 39618 28766
rect 39566 28690 39618 28702
rect 7646 28642 7698 28654
rect 5058 28590 5070 28642
rect 5122 28590 5134 28642
rect 7646 28578 7698 28590
rect 8878 28642 8930 28654
rect 8878 28578 8930 28590
rect 9102 28642 9154 28654
rect 9102 28578 9154 28590
rect 9326 28642 9378 28654
rect 9886 28642 9938 28654
rect 9538 28590 9550 28642
rect 9602 28590 9614 28642
rect 9326 28578 9378 28590
rect 9886 28578 9938 28590
rect 14590 28642 14642 28654
rect 14590 28578 14642 28590
rect 15150 28642 15202 28654
rect 15150 28578 15202 28590
rect 15486 28642 15538 28654
rect 16830 28642 16882 28654
rect 16370 28590 16382 28642
rect 16434 28590 16446 28642
rect 15486 28578 15538 28590
rect 16830 28578 16882 28590
rect 17838 28642 17890 28654
rect 26674 28590 26686 28642
rect 26738 28590 26750 28642
rect 29474 28590 29486 28642
rect 29538 28590 29550 28642
rect 17838 28578 17890 28590
rect 10446 28530 10498 28542
rect 34750 28530 34802 28542
rect 4274 28478 4286 28530
rect 4338 28478 4350 28530
rect 26898 28478 26910 28530
rect 26962 28478 26974 28530
rect 29698 28478 29710 28530
rect 29762 28478 29774 28530
rect 10446 28466 10498 28478
rect 34750 28466 34802 28478
rect 10110 28418 10162 28430
rect 10110 28354 10162 28366
rect 15934 28418 15986 28430
rect 15934 28354 15986 28366
rect 17390 28418 17442 28430
rect 17390 28354 17442 28366
rect 34974 28418 35026 28430
rect 34974 28354 35026 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 6302 28082 6354 28094
rect 6302 28018 6354 28030
rect 9438 28082 9490 28094
rect 9438 28018 9490 28030
rect 10782 28082 10834 28094
rect 10782 28018 10834 28030
rect 14030 28082 14082 28094
rect 14030 28018 14082 28030
rect 14142 28082 14194 28094
rect 14142 28018 14194 28030
rect 16606 28082 16658 28094
rect 22318 28082 22370 28094
rect 18162 28030 18174 28082
rect 18226 28030 18238 28082
rect 16606 28018 16658 28030
rect 22318 28018 22370 28030
rect 28590 28082 28642 28094
rect 28590 28018 28642 28030
rect 29150 28082 29202 28094
rect 29150 28018 29202 28030
rect 31278 28082 31330 28094
rect 31278 28018 31330 28030
rect 32398 28082 32450 28094
rect 32398 28018 32450 28030
rect 36318 28082 36370 28094
rect 36318 28018 36370 28030
rect 38782 28082 38834 28094
rect 38782 28018 38834 28030
rect 8094 27970 8146 27982
rect 5058 27918 5070 27970
rect 5122 27918 5134 27970
rect 8094 27906 8146 27918
rect 8990 27970 9042 27982
rect 8990 27906 9042 27918
rect 9550 27970 9602 27982
rect 9550 27906 9602 27918
rect 10446 27970 10498 27982
rect 20414 27970 20466 27982
rect 14242 27918 14254 27970
rect 14306 27918 14318 27970
rect 16370 27918 16382 27970
rect 16434 27918 16446 27970
rect 17938 27918 17950 27970
rect 18002 27918 18014 27970
rect 19842 27918 19854 27970
rect 19906 27918 19918 27970
rect 10446 27906 10498 27918
rect 20414 27906 20466 27918
rect 31502 27970 31554 27982
rect 31502 27906 31554 27918
rect 31614 27970 31666 27982
rect 31614 27906 31666 27918
rect 31838 27970 31890 27982
rect 31838 27906 31890 27918
rect 32174 27970 32226 27982
rect 39118 27970 39170 27982
rect 36642 27918 36654 27970
rect 36706 27918 36718 27970
rect 32174 27906 32226 27918
rect 39118 27906 39170 27918
rect 39342 27970 39394 27982
rect 39342 27906 39394 27918
rect 39902 27970 39954 27982
rect 39902 27906 39954 27918
rect 11342 27858 11394 27870
rect 15822 27858 15874 27870
rect 5730 27806 5742 27858
rect 5794 27806 5806 27858
rect 8754 27806 8766 27858
rect 8818 27806 8830 27858
rect 10210 27806 10222 27858
rect 10274 27806 10286 27858
rect 14802 27806 14814 27858
rect 14866 27806 14878 27858
rect 15026 27806 15038 27858
rect 15090 27806 15102 27858
rect 11342 27794 11394 27806
rect 15822 27794 15874 27806
rect 17502 27858 17554 27870
rect 20750 27858 20802 27870
rect 18386 27806 18398 27858
rect 18450 27806 18462 27858
rect 18834 27806 18846 27858
rect 18898 27806 18910 27858
rect 19282 27806 19294 27858
rect 19346 27806 19358 27858
rect 23090 27806 23102 27858
rect 23154 27806 23166 27858
rect 28130 27806 28142 27858
rect 28194 27806 28206 27858
rect 29362 27806 29374 27858
rect 29426 27806 29438 27858
rect 33058 27806 33070 27858
rect 33122 27806 33134 27858
rect 40226 27806 40238 27858
rect 40290 27806 40302 27858
rect 17502 27794 17554 27806
rect 20750 27794 20802 27806
rect 7646 27746 7698 27758
rect 2930 27694 2942 27746
rect 2994 27694 3006 27746
rect 7646 27682 7698 27694
rect 7758 27746 7810 27758
rect 7758 27682 7810 27694
rect 8206 27746 8258 27758
rect 8206 27682 8258 27694
rect 8318 27746 8370 27758
rect 8318 27682 8370 27694
rect 9774 27746 9826 27758
rect 9774 27682 9826 27694
rect 9998 27746 10050 27758
rect 9998 27682 10050 27694
rect 22766 27746 22818 27758
rect 22766 27682 22818 27694
rect 23886 27746 23938 27758
rect 23886 27682 23938 27694
rect 24782 27746 24834 27758
rect 29934 27746 29986 27758
rect 37102 27746 37154 27758
rect 25218 27694 25230 27746
rect 25282 27694 25294 27746
rect 27346 27694 27358 27746
rect 27410 27694 27422 27746
rect 32498 27694 32510 27746
rect 32562 27694 32574 27746
rect 33842 27694 33854 27746
rect 33906 27694 33918 27746
rect 35970 27694 35982 27746
rect 36034 27694 36046 27746
rect 24782 27682 24834 27694
rect 29934 27682 29986 27694
rect 37102 27682 37154 27694
rect 40014 27746 40066 27758
rect 40014 27682 40066 27694
rect 8542 27634 8594 27646
rect 23102 27634 23154 27646
rect 22306 27582 22318 27634
rect 22370 27631 22382 27634
rect 22754 27631 22766 27634
rect 22370 27585 22766 27631
rect 22370 27582 22382 27585
rect 22754 27582 22766 27585
rect 22818 27582 22830 27634
rect 8542 27570 8594 27582
rect 23102 27570 23154 27582
rect 23438 27634 23490 27646
rect 23438 27570 23490 27582
rect 39454 27634 39506 27646
rect 39454 27570 39506 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 6862 27298 6914 27310
rect 6862 27234 6914 27246
rect 21310 27298 21362 27310
rect 23998 27298 24050 27310
rect 26910 27298 26962 27310
rect 22306 27246 22318 27298
rect 22370 27246 22382 27298
rect 25890 27246 25902 27298
rect 25954 27246 25966 27298
rect 21310 27234 21362 27246
rect 23998 27234 24050 27246
rect 26910 27234 26962 27246
rect 5854 27186 5906 27198
rect 2146 27134 2158 27186
rect 2210 27134 2222 27186
rect 4274 27134 4286 27186
rect 4338 27134 4350 27186
rect 5854 27122 5906 27134
rect 9886 27186 9938 27198
rect 9886 27122 9938 27134
rect 11566 27186 11618 27198
rect 11566 27122 11618 27134
rect 19966 27186 20018 27198
rect 19966 27122 20018 27134
rect 21870 27186 21922 27198
rect 21870 27122 21922 27134
rect 26350 27186 26402 27198
rect 26350 27122 26402 27134
rect 27358 27186 27410 27198
rect 27358 27122 27410 27134
rect 31950 27186 32002 27198
rect 39778 27134 39790 27186
rect 39842 27134 39854 27186
rect 41906 27134 41918 27186
rect 41970 27134 41982 27186
rect 31950 27122 32002 27134
rect 10446 27074 10498 27086
rect 5058 27022 5070 27074
rect 5122 27022 5134 27074
rect 10446 27010 10498 27022
rect 11118 27074 11170 27086
rect 11118 27010 11170 27022
rect 14254 27074 14306 27086
rect 19406 27074 19458 27086
rect 14466 27022 14478 27074
rect 14530 27022 14542 27074
rect 15810 27022 15822 27074
rect 15874 27022 15886 27074
rect 16370 27022 16382 27074
rect 16434 27022 16446 27074
rect 17490 27022 17502 27074
rect 17554 27022 17566 27074
rect 18162 27022 18174 27074
rect 18226 27022 18238 27074
rect 18386 27022 18398 27074
rect 18450 27022 18462 27074
rect 14254 27010 14306 27022
rect 19406 27010 19458 27022
rect 20414 27074 20466 27086
rect 22878 27074 22930 27086
rect 21970 27022 21982 27074
rect 22034 27022 22046 27074
rect 22306 27022 22318 27074
rect 22370 27022 22382 27074
rect 20414 27010 20466 27022
rect 22878 27010 22930 27022
rect 23326 27074 23378 27086
rect 24110 27074 24162 27086
rect 25230 27074 25282 27086
rect 26462 27074 26514 27086
rect 23426 27022 23438 27074
rect 23490 27022 23502 27074
rect 24994 27022 25006 27074
rect 25058 27022 25070 27074
rect 25666 27022 25678 27074
rect 25730 27022 25742 27074
rect 26226 27022 26238 27074
rect 26290 27022 26302 27074
rect 23326 27010 23378 27022
rect 24110 27010 24162 27022
rect 25230 27010 25282 27022
rect 26462 27010 26514 27022
rect 35310 27074 35362 27086
rect 35310 27010 35362 27022
rect 35534 27074 35586 27086
rect 35534 27010 35586 27022
rect 36318 27074 36370 27086
rect 38994 27022 39006 27074
rect 39058 27022 39070 27074
rect 36318 27010 36370 27022
rect 6750 26962 6802 26974
rect 6750 26898 6802 26910
rect 10782 26962 10834 26974
rect 21422 26962 21474 26974
rect 15922 26910 15934 26962
rect 15986 26910 15998 26962
rect 16594 26910 16606 26962
rect 16658 26910 16670 26962
rect 17042 26910 17054 26962
rect 17106 26910 17118 26962
rect 19170 26910 19182 26962
rect 19234 26910 19246 26962
rect 10782 26898 10834 26910
rect 21422 26898 21474 26910
rect 21758 26962 21810 26974
rect 25342 26962 25394 26974
rect 23090 26910 23102 26962
rect 23154 26910 23166 26962
rect 21758 26898 21810 26910
rect 25342 26898 25394 26910
rect 26798 26962 26850 26974
rect 26798 26898 26850 26910
rect 35870 26962 35922 26974
rect 35870 26898 35922 26910
rect 14366 26850 14418 26862
rect 14366 26786 14418 26798
rect 16942 26850 16994 26862
rect 16942 26786 16994 26798
rect 23662 26850 23714 26862
rect 23662 26786 23714 26798
rect 24222 26850 24274 26862
rect 24222 26786 24274 26798
rect 35758 26850 35810 26862
rect 35758 26786 35810 26798
rect 38670 26850 38722 26862
rect 38670 26786 38722 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 17614 26514 17666 26526
rect 17614 26450 17666 26462
rect 19406 26514 19458 26526
rect 22542 26514 22594 26526
rect 36206 26514 36258 26526
rect 19842 26462 19854 26514
rect 19906 26462 19918 26514
rect 23314 26462 23326 26514
rect 23378 26462 23390 26514
rect 19406 26450 19458 26462
rect 22542 26450 22594 26462
rect 36206 26450 36258 26462
rect 7982 26402 8034 26414
rect 7982 26338 8034 26350
rect 8878 26402 8930 26414
rect 16270 26402 16322 26414
rect 36766 26402 36818 26414
rect 9762 26350 9774 26402
rect 9826 26350 9838 26402
rect 19618 26350 19630 26402
rect 19682 26350 19694 26402
rect 21522 26350 21534 26402
rect 21586 26350 21598 26402
rect 8878 26338 8930 26350
rect 16270 26338 16322 26350
rect 36766 26338 36818 26350
rect 8430 26290 8482 26302
rect 15262 26290 15314 26302
rect 4050 26238 4062 26290
rect 4114 26238 4126 26290
rect 8642 26238 8654 26290
rect 8706 26238 8718 26290
rect 9986 26238 9998 26290
rect 10050 26238 10062 26290
rect 8430 26226 8482 26238
rect 15262 26226 15314 26238
rect 15822 26290 15874 26302
rect 21198 26290 21250 26302
rect 19954 26238 19966 26290
rect 20018 26238 20030 26290
rect 20738 26238 20750 26290
rect 20802 26238 20814 26290
rect 15822 26226 15874 26238
rect 21198 26226 21250 26238
rect 21982 26290 22034 26302
rect 21982 26226 22034 26238
rect 22878 26290 22930 26302
rect 36542 26290 36594 26302
rect 23090 26238 23102 26290
rect 23154 26238 23166 26290
rect 23650 26238 23662 26290
rect 23714 26238 23726 26290
rect 24322 26238 24334 26290
rect 24386 26238 24398 26290
rect 37202 26238 37214 26290
rect 37266 26238 37278 26290
rect 22878 26226 22930 26238
rect 36542 26226 36594 26238
rect 1934 26178 1986 26190
rect 1934 26114 1986 26126
rect 8094 26178 8146 26190
rect 8094 26114 8146 26126
rect 8206 26178 8258 26190
rect 8206 26114 8258 26126
rect 16718 26178 16770 26190
rect 16718 26114 16770 26126
rect 24110 26178 24162 26190
rect 24110 26114 24162 26126
rect 25342 26178 25394 26190
rect 25342 26114 25394 26126
rect 33182 26178 33234 26190
rect 33182 26114 33234 26126
rect 33742 26178 33794 26190
rect 36866 26126 36878 26178
rect 36930 26126 36942 26178
rect 37986 26126 37998 26178
rect 38050 26126 38062 26178
rect 40226 26126 40238 26178
rect 40290 26126 40302 26178
rect 33742 26114 33794 26126
rect 23998 26066 24050 26078
rect 23426 26014 23438 26066
rect 23490 26014 23502 26066
rect 23998 26002 24050 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 6862 25730 6914 25742
rect 6862 25666 6914 25678
rect 33518 25730 33570 25742
rect 33518 25666 33570 25678
rect 34526 25730 34578 25742
rect 34526 25666 34578 25678
rect 1934 25618 1986 25630
rect 1934 25554 1986 25566
rect 14926 25618 14978 25630
rect 16494 25618 16546 25630
rect 32846 25618 32898 25630
rect 15698 25566 15710 25618
rect 15762 25566 15774 25618
rect 23202 25566 23214 25618
rect 23266 25566 23278 25618
rect 29474 25566 29486 25618
rect 29538 25566 29550 25618
rect 14926 25554 14978 25566
rect 16494 25554 16546 25566
rect 32846 25554 32898 25566
rect 35758 25618 35810 25630
rect 35758 25554 35810 25566
rect 14702 25506 14754 25518
rect 34638 25506 34690 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 14018 25454 14030 25506
rect 14082 25454 14094 25506
rect 17602 25454 17614 25506
rect 17666 25454 17678 25506
rect 18946 25454 18958 25506
rect 19010 25454 19022 25506
rect 19506 25454 19518 25506
rect 19570 25454 19582 25506
rect 20402 25454 20414 25506
rect 20466 25454 20478 25506
rect 26786 25454 26798 25506
rect 26850 25454 26862 25506
rect 32386 25454 32398 25506
rect 32450 25454 32462 25506
rect 33394 25454 33406 25506
rect 33458 25454 33470 25506
rect 33618 25454 33630 25506
rect 33682 25454 33694 25506
rect 33954 25454 33966 25506
rect 34018 25454 34030 25506
rect 14702 25442 14754 25454
rect 34638 25442 34690 25454
rect 35086 25506 35138 25518
rect 35086 25442 35138 25454
rect 35310 25506 35362 25518
rect 35310 25442 35362 25454
rect 38894 25506 38946 25518
rect 38894 25442 38946 25454
rect 39342 25506 39394 25518
rect 39342 25442 39394 25454
rect 39566 25506 39618 25518
rect 39566 25442 39618 25454
rect 40126 25506 40178 25518
rect 40126 25442 40178 25454
rect 6750 25394 6802 25406
rect 14814 25394 14866 25406
rect 14242 25342 14254 25394
rect 14306 25342 14318 25394
rect 6750 25330 6802 25342
rect 14814 25330 14866 25342
rect 15038 25394 15090 25406
rect 15038 25330 15090 25342
rect 15934 25394 15986 25406
rect 34190 25394 34242 25406
rect 17714 25342 17726 25394
rect 17778 25342 17790 25394
rect 19730 25342 19742 25394
rect 19794 25342 19806 25394
rect 20290 25342 20302 25394
rect 20354 25342 20366 25394
rect 31602 25342 31614 25394
rect 31666 25342 31678 25394
rect 15934 25330 15986 25342
rect 34190 25330 34242 25342
rect 34414 25394 34466 25406
rect 34414 25330 34466 25342
rect 34862 25394 34914 25406
rect 34862 25330 34914 25342
rect 47854 25394 47906 25406
rect 47854 25330 47906 25342
rect 48190 25394 48242 25406
rect 48190 25330 48242 25342
rect 15150 25282 15202 25294
rect 15150 25218 15202 25230
rect 15710 25282 15762 25294
rect 15710 25218 15762 25230
rect 17166 25282 17218 25294
rect 18398 25282 18450 25294
rect 17826 25230 17838 25282
rect 17890 25230 17902 25282
rect 17166 25218 17218 25230
rect 18398 25218 18450 25230
rect 27246 25282 27298 25294
rect 27246 25218 27298 25230
rect 33182 25282 33234 25294
rect 33182 25218 33234 25230
rect 39118 25282 39170 25294
rect 39118 25218 39170 25230
rect 47630 25282 47682 25294
rect 47630 25218 47682 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 16494 24946 16546 24958
rect 14802 24894 14814 24946
rect 14866 24894 14878 24946
rect 16494 24882 16546 24894
rect 16606 24946 16658 24958
rect 16606 24882 16658 24894
rect 17614 24946 17666 24958
rect 17614 24882 17666 24894
rect 18510 24946 18562 24958
rect 18510 24882 18562 24894
rect 22318 24946 22370 24958
rect 22318 24882 22370 24894
rect 33294 24946 33346 24958
rect 33294 24882 33346 24894
rect 34638 24946 34690 24958
rect 34638 24882 34690 24894
rect 34974 24946 35026 24958
rect 34974 24882 35026 24894
rect 13358 24834 13410 24846
rect 4946 24782 4958 24834
rect 5010 24782 5022 24834
rect 11666 24782 11678 24834
rect 11730 24782 11742 24834
rect 13358 24770 13410 24782
rect 19854 24834 19906 24846
rect 34862 24834 34914 24846
rect 23986 24782 23998 24834
rect 24050 24782 24062 24834
rect 19854 24770 19906 24782
rect 34862 24770 34914 24782
rect 36318 24834 36370 24846
rect 39678 24834 39730 24846
rect 39106 24782 39118 24834
rect 39170 24831 39182 24834
rect 39330 24831 39342 24834
rect 39170 24785 39342 24831
rect 39170 24782 39182 24785
rect 39330 24782 39342 24785
rect 39394 24782 39406 24834
rect 36318 24770 36370 24782
rect 39678 24770 39730 24782
rect 16046 24722 16098 24734
rect 16718 24722 16770 24734
rect 5730 24670 5742 24722
rect 5794 24670 5806 24722
rect 11778 24670 11790 24722
rect 11842 24670 11854 24722
rect 12450 24670 12462 24722
rect 12514 24670 12526 24722
rect 12786 24670 12798 24722
rect 12850 24670 12862 24722
rect 16370 24670 16382 24722
rect 16434 24670 16446 24722
rect 16046 24658 16098 24670
rect 16718 24658 16770 24670
rect 17950 24722 18002 24734
rect 18398 24722 18450 24734
rect 18274 24670 18286 24722
rect 18338 24670 18350 24722
rect 17950 24658 18002 24670
rect 18398 24658 18450 24670
rect 18622 24722 18674 24734
rect 31054 24722 31106 24734
rect 23762 24670 23774 24722
rect 23826 24670 23838 24722
rect 30482 24670 30494 24722
rect 30546 24670 30558 24722
rect 18622 24658 18674 24670
rect 31054 24658 31106 24670
rect 33630 24722 33682 24734
rect 33630 24658 33682 24670
rect 34302 24722 34354 24734
rect 39454 24722 39506 24734
rect 36642 24670 36654 24722
rect 36706 24670 36718 24722
rect 34302 24658 34354 24670
rect 39454 24658 39506 24670
rect 6302 24610 6354 24622
rect 14590 24610 14642 24622
rect 2818 24558 2830 24610
rect 2882 24558 2894 24610
rect 11890 24558 11902 24610
rect 11954 24558 11966 24610
rect 6302 24546 6354 24558
rect 14590 24546 14642 24558
rect 19182 24610 19234 24622
rect 34078 24610 34130 24622
rect 20290 24558 20302 24610
rect 20354 24558 20366 24610
rect 27570 24558 27582 24610
rect 27634 24558 27646 24610
rect 29698 24558 29710 24610
rect 29762 24558 29774 24610
rect 19182 24546 19234 24558
rect 34078 24546 34130 24558
rect 36654 24498 36706 24510
rect 36654 24434 36706 24446
rect 39790 24498 39842 24510
rect 39790 24434 39842 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 13022 24162 13074 24174
rect 13022 24098 13074 24110
rect 23774 24162 23826 24174
rect 23774 24098 23826 24110
rect 1934 24050 1986 24062
rect 1934 23986 1986 23998
rect 7646 24050 7698 24062
rect 7646 23986 7698 23998
rect 28590 24050 28642 24062
rect 28590 23986 28642 23998
rect 29822 24050 29874 24062
rect 29822 23986 29874 23998
rect 34078 24050 34130 24062
rect 34078 23986 34130 23998
rect 36430 24050 36482 24062
rect 39902 24050 39954 24062
rect 43374 24050 43426 24062
rect 37762 23998 37774 24050
rect 37826 23998 37838 24050
rect 41234 23998 41246 24050
rect 41298 23998 41310 24050
rect 36430 23986 36482 23998
rect 39902 23986 39954 23998
rect 43374 23986 43426 23998
rect 7198 23938 7250 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 7198 23874 7250 23886
rect 7422 23938 7474 23950
rect 8206 23938 8258 23950
rect 29486 23938 29538 23950
rect 7858 23886 7870 23938
rect 7922 23886 7934 23938
rect 11554 23886 11566 23938
rect 11618 23886 11630 23938
rect 12226 23886 12238 23938
rect 12290 23886 12302 23938
rect 12786 23886 12798 23938
rect 12850 23886 12862 23938
rect 13906 23886 13918 23938
rect 13970 23886 13982 23938
rect 17714 23886 17726 23938
rect 17778 23886 17790 23938
rect 25106 23886 25118 23938
rect 25170 23886 25182 23938
rect 29138 23886 29150 23938
rect 29202 23886 29214 23938
rect 7422 23874 7474 23886
rect 8206 23874 8258 23886
rect 29486 23874 29538 23886
rect 29598 23938 29650 23950
rect 30718 23938 30770 23950
rect 31502 23938 31554 23950
rect 30482 23886 30494 23938
rect 30546 23886 30558 23938
rect 30818 23886 30830 23938
rect 30882 23886 30894 23938
rect 37090 23886 37102 23938
rect 37154 23886 37166 23938
rect 40450 23886 40462 23938
rect 40514 23886 40526 23938
rect 29598 23874 29650 23886
rect 30718 23874 30770 23886
rect 31502 23874 31554 23886
rect 16494 23826 16546 23838
rect 12674 23774 12686 23826
rect 12738 23774 12750 23826
rect 14018 23774 14030 23826
rect 14082 23774 14094 23826
rect 16494 23762 16546 23774
rect 23326 23826 23378 23838
rect 23326 23762 23378 23774
rect 23662 23826 23714 23838
rect 23662 23762 23714 23774
rect 23774 23826 23826 23838
rect 23774 23762 23826 23774
rect 24222 23826 24274 23838
rect 24222 23762 24274 23774
rect 24558 23826 24610 23838
rect 24558 23762 24610 23774
rect 24894 23826 24946 23838
rect 24894 23762 24946 23774
rect 29934 23826 29986 23838
rect 29934 23762 29986 23774
rect 30270 23826 30322 23838
rect 30270 23762 30322 23774
rect 7646 23714 7698 23726
rect 7646 23650 7698 23662
rect 8542 23714 8594 23726
rect 31054 23714 31106 23726
rect 15474 23662 15486 23714
rect 15538 23662 15550 23714
rect 8542 23650 8594 23662
rect 31054 23650 31106 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 24670 23378 24722 23390
rect 24670 23314 24722 23326
rect 27582 23378 27634 23390
rect 27582 23314 27634 23326
rect 40126 23378 40178 23390
rect 40126 23314 40178 23326
rect 5742 23266 5794 23278
rect 5742 23202 5794 23214
rect 7086 23266 7138 23278
rect 15262 23266 15314 23278
rect 27694 23266 27746 23278
rect 12674 23214 12686 23266
rect 12738 23214 12750 23266
rect 17378 23214 17390 23266
rect 17442 23214 17454 23266
rect 20402 23214 20414 23266
rect 20466 23214 20478 23266
rect 25554 23214 25566 23266
rect 25618 23214 25630 23266
rect 7086 23202 7138 23214
rect 15262 23202 15314 23214
rect 27694 23202 27746 23214
rect 30270 23266 30322 23278
rect 30270 23202 30322 23214
rect 5854 23154 5906 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 5854 23090 5906 23102
rect 7310 23154 7362 23166
rect 7310 23090 7362 23102
rect 7534 23154 7586 23166
rect 8878 23154 8930 23166
rect 7746 23102 7758 23154
rect 7810 23102 7822 23154
rect 7970 23102 7982 23154
rect 8034 23102 8046 23154
rect 7534 23090 7586 23102
rect 8878 23090 8930 23102
rect 11678 23154 11730 23166
rect 14702 23154 14754 23166
rect 21198 23154 21250 23166
rect 27134 23154 27186 23166
rect 12562 23102 12574 23154
rect 12626 23102 12638 23154
rect 17490 23102 17502 23154
rect 17554 23102 17566 23154
rect 18162 23102 18174 23154
rect 18226 23102 18238 23154
rect 18610 23102 18622 23154
rect 18674 23102 18686 23154
rect 20290 23102 20302 23154
rect 20354 23102 20366 23154
rect 25218 23102 25230 23154
rect 25282 23102 25294 23154
rect 28242 23102 28254 23154
rect 28306 23102 28318 23154
rect 11678 23090 11730 23102
rect 14702 23090 14754 23102
rect 21198 23090 21250 23102
rect 27134 23090 27186 23102
rect 5182 23042 5234 23054
rect 5182 22978 5234 22990
rect 7198 23042 7250 23054
rect 8654 23042 8706 23054
rect 8306 22990 8318 23042
rect 8370 22990 8382 23042
rect 7198 22978 7250 22990
rect 8654 22978 8706 22990
rect 9774 23042 9826 23054
rect 9774 22978 9826 22990
rect 12238 23042 12290 23054
rect 28702 23042 28754 23054
rect 13794 22990 13806 23042
rect 13858 22990 13870 23042
rect 20738 22990 20750 23042
rect 20802 22990 20814 23042
rect 25778 22990 25790 23042
rect 25842 22990 25854 23042
rect 12238 22978 12290 22990
rect 28702 22978 28754 22990
rect 29710 23042 29762 23054
rect 30370 22990 30382 23042
rect 30434 22990 30446 23042
rect 29710 22978 29762 22990
rect 1934 22930 1986 22942
rect 27470 22930 27522 22942
rect 18498 22878 18510 22930
rect 18562 22878 18574 22930
rect 1934 22866 1986 22878
rect 27470 22866 27522 22878
rect 30046 22930 30098 22942
rect 30046 22866 30098 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 5966 22594 6018 22606
rect 5966 22530 6018 22542
rect 9886 22482 9938 22494
rect 2034 22430 2046 22482
rect 2098 22430 2110 22482
rect 4162 22430 4174 22482
rect 4226 22430 4238 22482
rect 9886 22418 9938 22430
rect 11118 22482 11170 22494
rect 14366 22482 14418 22494
rect 12002 22430 12014 22482
rect 12066 22430 12078 22482
rect 11118 22418 11170 22430
rect 14366 22418 14418 22430
rect 16382 22482 16434 22494
rect 18622 22482 18674 22494
rect 23774 22482 23826 22494
rect 18274 22430 18286 22482
rect 18338 22430 18350 22482
rect 21746 22430 21758 22482
rect 21810 22430 21822 22482
rect 16382 22418 16434 22430
rect 18622 22418 18674 22430
rect 23774 22418 23826 22430
rect 8990 22370 9042 22382
rect 14030 22370 14082 22382
rect 4946 22318 4958 22370
rect 5010 22318 5022 22370
rect 10658 22318 10670 22370
rect 10722 22318 10734 22370
rect 12562 22318 12574 22370
rect 12626 22318 12638 22370
rect 8990 22306 9042 22318
rect 14030 22306 14082 22318
rect 16046 22370 16098 22382
rect 29586 22318 29598 22370
rect 29650 22318 29662 22370
rect 16046 22306 16098 22318
rect 5854 22258 5906 22270
rect 5854 22194 5906 22206
rect 8766 22258 8818 22270
rect 8766 22194 8818 22206
rect 13582 22258 13634 22270
rect 13582 22194 13634 22206
rect 14254 22258 14306 22270
rect 14254 22194 14306 22206
rect 15150 22258 15202 22270
rect 15150 22194 15202 22206
rect 18398 22258 18450 22270
rect 24670 22258 24722 22270
rect 23426 22206 23438 22258
rect 23490 22206 23502 22258
rect 18398 22194 18450 22206
rect 24670 22194 24722 22206
rect 25230 22258 25282 22270
rect 25230 22194 25282 22206
rect 8318 22146 8370 22158
rect 8318 22082 8370 22094
rect 9102 22146 9154 22158
rect 9102 22082 9154 22094
rect 9214 22146 9266 22158
rect 9214 22082 9266 22094
rect 9326 22146 9378 22158
rect 9326 22082 9378 22094
rect 13806 22146 13858 22158
rect 20862 22146 20914 22158
rect 16594 22094 16606 22146
rect 16658 22094 16670 22146
rect 13806 22082 13858 22094
rect 20862 22082 20914 22094
rect 21310 22146 21362 22158
rect 21310 22082 21362 22094
rect 23102 22146 23154 22158
rect 23102 22082 23154 22094
rect 24334 22146 24386 22158
rect 24334 22082 24386 22094
rect 24782 22146 24834 22158
rect 24782 22082 24834 22094
rect 25006 22146 25058 22158
rect 25006 22082 25058 22094
rect 25342 22146 25394 22158
rect 25342 22082 25394 22094
rect 25566 22146 25618 22158
rect 25566 22082 25618 22094
rect 25902 22146 25954 22158
rect 29810 22094 29822 22146
rect 29874 22094 29886 22146
rect 25902 22082 25954 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 16606 21810 16658 21822
rect 11442 21758 11454 21810
rect 11506 21758 11518 21810
rect 16606 21746 16658 21758
rect 19630 21810 19682 21822
rect 24670 21810 24722 21822
rect 22194 21758 22206 21810
rect 22258 21758 22270 21810
rect 23874 21758 23886 21810
rect 23938 21758 23950 21810
rect 19630 21746 19682 21758
rect 24670 21746 24722 21758
rect 34414 21810 34466 21822
rect 34414 21746 34466 21758
rect 35198 21810 35250 21822
rect 35198 21746 35250 21758
rect 37886 21810 37938 21822
rect 37886 21746 37938 21758
rect 8990 21698 9042 21710
rect 12574 21698 12626 21710
rect 10098 21646 10110 21698
rect 10162 21646 10174 21698
rect 8990 21634 9042 21646
rect 12574 21634 12626 21646
rect 15710 21698 15762 21710
rect 15710 21634 15762 21646
rect 19854 21698 19906 21710
rect 21534 21698 21586 21710
rect 20738 21646 20750 21698
rect 20802 21646 20814 21698
rect 19854 21634 19906 21646
rect 21534 21634 21586 21646
rect 22878 21698 22930 21710
rect 34738 21646 34750 21698
rect 34802 21646 34814 21698
rect 22878 21634 22930 21646
rect 8430 21586 8482 21598
rect 4386 21534 4398 21586
rect 4450 21534 4462 21586
rect 5170 21534 5182 21586
rect 5234 21534 5246 21586
rect 8430 21522 8482 21534
rect 9550 21586 9602 21598
rect 9550 21522 9602 21534
rect 9662 21586 9714 21598
rect 12126 21586 12178 21598
rect 11554 21534 11566 21586
rect 11618 21534 11630 21586
rect 9662 21522 9714 21534
rect 12126 21522 12178 21534
rect 16606 21586 16658 21598
rect 16606 21522 16658 21534
rect 19406 21586 19458 21598
rect 19406 21522 19458 21534
rect 19966 21586 20018 21598
rect 19966 21522 20018 21534
rect 21086 21586 21138 21598
rect 21086 21522 21138 21534
rect 21310 21586 21362 21598
rect 21310 21522 21362 21534
rect 21646 21586 21698 21598
rect 21646 21522 21698 21534
rect 22542 21586 22594 21598
rect 22542 21522 22594 21534
rect 23214 21586 23266 21598
rect 23650 21534 23662 21586
rect 23714 21534 23726 21586
rect 23214 21522 23266 21534
rect 5630 21474 5682 21486
rect 2258 21422 2270 21474
rect 2322 21422 2334 21474
rect 5630 21410 5682 21422
rect 7646 21474 7698 21486
rect 7646 21410 7698 21422
rect 8094 21474 8146 21486
rect 8094 21410 8146 21422
rect 14926 21474 14978 21486
rect 14926 21410 14978 21422
rect 20526 21474 20578 21486
rect 20526 21410 20578 21422
rect 25342 21474 25394 21486
rect 25342 21410 25394 21422
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 12898 20974 12910 21026
rect 12962 20974 12974 21026
rect 22866 20974 22878 21026
rect 22930 20974 22942 21026
rect 1934 20914 1986 20926
rect 1934 20850 1986 20862
rect 9998 20914 10050 20926
rect 9998 20850 10050 20862
rect 10894 20914 10946 20926
rect 10894 20850 10946 20862
rect 12014 20914 12066 20926
rect 12014 20850 12066 20862
rect 12350 20914 12402 20926
rect 21534 20914 21586 20926
rect 18050 20862 18062 20914
rect 18114 20862 18126 20914
rect 12350 20850 12402 20862
rect 21534 20850 21586 20862
rect 24558 20914 24610 20926
rect 24558 20850 24610 20862
rect 25566 20914 25618 20926
rect 34974 20914 35026 20926
rect 30930 20862 30942 20914
rect 30994 20862 31006 20914
rect 25566 20850 25618 20862
rect 34974 20850 35026 20862
rect 41134 20914 41186 20926
rect 41134 20850 41186 20862
rect 10334 20802 10386 20814
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 10334 20738 10386 20750
rect 12574 20802 12626 20814
rect 12574 20738 12626 20750
rect 14366 20802 14418 20814
rect 22318 20802 22370 20814
rect 15362 20750 15374 20802
rect 15426 20750 15438 20802
rect 17938 20750 17950 20802
rect 18002 20750 18014 20802
rect 14366 20738 14418 20750
rect 22318 20738 22370 20750
rect 22542 20802 22594 20814
rect 22542 20738 22594 20750
rect 23774 20802 23826 20814
rect 23774 20738 23826 20750
rect 25342 20802 25394 20814
rect 25342 20738 25394 20750
rect 29374 20802 29426 20814
rect 29374 20738 29426 20750
rect 29934 20802 29986 20814
rect 34190 20802 34242 20814
rect 37550 20802 37602 20814
rect 33842 20750 33854 20802
rect 33906 20750 33918 20802
rect 35522 20750 35534 20802
rect 35586 20750 35598 20802
rect 38210 20750 38222 20802
rect 38274 20750 38286 20802
rect 29934 20738 29986 20750
rect 34190 20738 34242 20750
rect 37550 20738 37602 20750
rect 20414 20690 20466 20702
rect 15586 20638 15598 20690
rect 15650 20638 15662 20690
rect 16258 20638 16270 20690
rect 16322 20638 16334 20690
rect 30158 20690 30210 20702
rect 20414 20626 20466 20638
rect 29710 20634 29762 20646
rect 9102 20578 9154 20590
rect 9102 20514 9154 20526
rect 9438 20578 9490 20590
rect 9438 20514 9490 20526
rect 11454 20578 11506 20590
rect 11454 20514 11506 20526
rect 13806 20578 13858 20590
rect 13806 20514 13858 20526
rect 21982 20578 22034 20590
rect 21982 20514 22034 20526
rect 23214 20578 23266 20590
rect 23214 20514 23266 20526
rect 25006 20578 25058 20590
rect 28590 20578 28642 20590
rect 25890 20526 25902 20578
rect 25954 20526 25966 20578
rect 25006 20514 25058 20526
rect 28590 20514 28642 20526
rect 29598 20578 29650 20590
rect 30158 20626 30210 20638
rect 30382 20690 30434 20702
rect 30382 20626 30434 20638
rect 30606 20690 30658 20702
rect 36990 20690 37042 20702
rect 33058 20638 33070 20690
rect 33122 20638 33134 20690
rect 30606 20626 30658 20638
rect 36990 20626 37042 20638
rect 37214 20690 37266 20702
rect 37214 20626 37266 20638
rect 37438 20690 37490 20702
rect 38994 20638 39006 20690
rect 39058 20638 39070 20690
rect 37438 20626 37490 20638
rect 29710 20570 29762 20582
rect 35758 20578 35810 20590
rect 34514 20526 34526 20578
rect 34578 20526 34590 20578
rect 29598 20514 29650 20526
rect 35758 20514 35810 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 12238 20242 12290 20254
rect 12238 20178 12290 20190
rect 24222 20242 24274 20254
rect 24222 20178 24274 20190
rect 30494 20242 30546 20254
rect 30494 20178 30546 20190
rect 2046 20130 2098 20142
rect 10110 20130 10162 20142
rect 8978 20078 8990 20130
rect 9042 20078 9054 20130
rect 2046 20066 2098 20078
rect 10110 20066 10162 20078
rect 11678 20130 11730 20142
rect 15374 20130 15426 20142
rect 12898 20078 12910 20130
rect 12962 20078 12974 20130
rect 14690 20078 14702 20130
rect 14754 20078 14766 20130
rect 11678 20066 11730 20078
rect 15374 20066 15426 20078
rect 24670 20130 24722 20142
rect 24670 20066 24722 20078
rect 26350 20130 26402 20142
rect 26350 20066 26402 20078
rect 26462 20130 26514 20142
rect 26462 20066 26514 20078
rect 27022 20130 27074 20142
rect 27022 20066 27074 20078
rect 30718 20130 30770 20142
rect 30718 20066 30770 20078
rect 31838 20130 31890 20142
rect 31838 20066 31890 20078
rect 34526 20130 34578 20142
rect 34526 20066 34578 20078
rect 34974 20130 35026 20142
rect 34974 20066 35026 20078
rect 35534 20130 35586 20142
rect 35534 20066 35586 20078
rect 35758 20130 35810 20142
rect 35758 20066 35810 20078
rect 47854 20130 47906 20142
rect 47854 20066 47906 20078
rect 1710 20018 1762 20030
rect 20750 20018 20802 20030
rect 8754 19966 8766 20018
rect 8818 19966 8830 20018
rect 12786 19966 12798 20018
rect 12850 19966 12862 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 1710 19954 1762 19966
rect 20750 19954 20802 19966
rect 21310 20018 21362 20030
rect 21310 19954 21362 19966
rect 25454 20018 25506 20030
rect 25454 19954 25506 19966
rect 25678 20018 25730 20030
rect 25678 19954 25730 19966
rect 26686 20018 26738 20030
rect 26686 19954 26738 19966
rect 30830 20018 30882 20030
rect 34862 20018 34914 20030
rect 32050 19966 32062 20018
rect 32114 19966 32126 20018
rect 30830 19954 30882 19966
rect 34862 19954 34914 19966
rect 35198 20018 35250 20030
rect 35198 19954 35250 19966
rect 35422 20018 35474 20030
rect 35422 19954 35474 19966
rect 36318 20018 36370 20030
rect 36318 19954 36370 19966
rect 36542 20018 36594 20030
rect 36542 19954 36594 19966
rect 36766 20018 36818 20030
rect 48190 20018 48242 20030
rect 37314 19966 37326 20018
rect 37378 19966 37390 20018
rect 36766 19954 36818 19966
rect 48190 19954 48242 19966
rect 2494 19906 2546 19918
rect 2494 19842 2546 19854
rect 7982 19906 8034 19918
rect 7982 19842 8034 19854
rect 8318 19906 8370 19918
rect 8318 19842 8370 19854
rect 9774 19906 9826 19918
rect 9774 19842 9826 19854
rect 10670 19906 10722 19918
rect 10670 19842 10722 19854
rect 11006 19906 11058 19918
rect 11902 19906 11954 19918
rect 11330 19854 11342 19906
rect 11394 19854 11406 19906
rect 11006 19842 11058 19854
rect 11902 19842 11954 19854
rect 20414 19906 20466 19918
rect 20414 19842 20466 19854
rect 22878 19906 22930 19918
rect 22878 19842 22930 19854
rect 23326 19906 23378 19918
rect 23326 19842 23378 19854
rect 30270 19906 30322 19918
rect 30270 19842 30322 19854
rect 36430 19906 36482 19918
rect 40126 19906 40178 19918
rect 37986 19854 37998 19906
rect 38050 19854 38062 19906
rect 36430 19842 36482 19854
rect 40126 19842 40178 19854
rect 47630 19906 47682 19918
rect 47630 19842 47682 19854
rect 22866 19742 22878 19794
rect 22930 19791 22942 19794
rect 23202 19791 23214 19794
rect 22930 19745 23214 19791
rect 22930 19742 22942 19745
rect 23202 19742 23214 19745
rect 23266 19742 23278 19794
rect 26002 19742 26014 19794
rect 26066 19742 26078 19794
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 12462 19458 12514 19470
rect 11554 19406 11566 19458
rect 11618 19406 11630 19458
rect 12462 19394 12514 19406
rect 14030 19458 14082 19470
rect 15934 19458 15986 19470
rect 14354 19406 14366 19458
rect 14418 19406 14430 19458
rect 14030 19394 14082 19406
rect 15934 19394 15986 19406
rect 36318 19458 36370 19470
rect 36318 19394 36370 19406
rect 37102 19458 37154 19470
rect 37102 19394 37154 19406
rect 10670 19346 10722 19358
rect 10670 19282 10722 19294
rect 12350 19346 12402 19358
rect 12350 19282 12402 19294
rect 13806 19346 13858 19358
rect 13806 19282 13858 19294
rect 16158 19346 16210 19358
rect 16158 19282 16210 19294
rect 16718 19346 16770 19358
rect 16718 19282 16770 19294
rect 19966 19346 20018 19358
rect 19966 19282 20018 19294
rect 27918 19346 27970 19358
rect 27918 19282 27970 19294
rect 35198 19346 35250 19358
rect 35198 19282 35250 19294
rect 37662 19346 37714 19358
rect 37662 19282 37714 19294
rect 38110 19346 38162 19358
rect 38110 19282 38162 19294
rect 9774 19234 9826 19246
rect 12014 19234 12066 19246
rect 10994 19182 11006 19234
rect 11058 19182 11070 19234
rect 9774 19170 9826 19182
rect 12014 19170 12066 19182
rect 12126 19234 12178 19246
rect 12126 19170 12178 19182
rect 15262 19234 15314 19246
rect 15262 19170 15314 19182
rect 26798 19234 26850 19246
rect 26798 19170 26850 19182
rect 30606 19234 30658 19246
rect 36430 19234 36482 19246
rect 31938 19182 31950 19234
rect 32002 19182 32014 19234
rect 30606 19170 30658 19182
rect 36430 19170 36482 19182
rect 36990 19234 37042 19246
rect 36990 19170 37042 19182
rect 15150 19122 15202 19134
rect 15150 19058 15202 19070
rect 19406 19122 19458 19134
rect 19406 19058 19458 19070
rect 19518 19122 19570 19134
rect 19518 19058 19570 19070
rect 27246 19122 27298 19134
rect 27246 19058 27298 19070
rect 27470 19122 27522 19134
rect 27470 19058 27522 19070
rect 31278 19122 31330 19134
rect 37102 19122 37154 19134
rect 31714 19070 31726 19122
rect 31778 19070 31790 19122
rect 31278 19058 31330 19070
rect 37102 19058 37154 19070
rect 8878 19010 8930 19022
rect 8878 18946 8930 18958
rect 9214 19010 9266 19022
rect 9214 18946 9266 18958
rect 10110 19010 10162 19022
rect 10110 18946 10162 18958
rect 14926 19010 14978 19022
rect 18174 19010 18226 19022
rect 15586 18958 15598 19010
rect 15650 18958 15662 19010
rect 14926 18946 14978 18958
rect 18174 18946 18226 18958
rect 19182 19010 19234 19022
rect 19182 18946 19234 18958
rect 27134 19010 27186 19022
rect 27134 18946 27186 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 30718 19010 30770 19022
rect 30718 18946 30770 18958
rect 30942 19010 30994 19022
rect 30942 18946 30994 18958
rect 32734 19010 32786 19022
rect 32734 18946 32786 18958
rect 35870 19010 35922 19022
rect 35870 18946 35922 18958
rect 36318 19010 36370 19022
rect 36318 18946 36370 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 11118 18674 11170 18686
rect 11118 18610 11170 18622
rect 15150 18674 15202 18686
rect 15150 18610 15202 18622
rect 16270 18674 16322 18686
rect 25666 18622 25678 18674
rect 25730 18622 25742 18674
rect 16270 18610 16322 18622
rect 2046 18562 2098 18574
rect 2046 18498 2098 18510
rect 9774 18562 9826 18574
rect 9774 18498 9826 18510
rect 11566 18562 11618 18574
rect 11566 18498 11618 18510
rect 13022 18562 13074 18574
rect 18062 18562 18114 18574
rect 15586 18510 15598 18562
rect 15650 18510 15662 18562
rect 13022 18498 13074 18510
rect 18062 18498 18114 18510
rect 18174 18562 18226 18574
rect 27906 18510 27918 18562
rect 27970 18510 27982 18562
rect 29362 18510 29374 18562
rect 29426 18510 29438 18562
rect 37650 18510 37662 18562
rect 37714 18510 37726 18562
rect 18174 18498 18226 18510
rect 1710 18450 1762 18462
rect 7198 18450 7250 18462
rect 24110 18450 24162 18462
rect 29038 18450 29090 18462
rect 6514 18398 6526 18450
rect 6578 18398 6590 18450
rect 11890 18398 11902 18450
rect 11954 18398 11966 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 28690 18398 28702 18450
rect 28754 18398 28766 18450
rect 1710 18386 1762 18398
rect 7198 18386 7250 18398
rect 24110 18386 24162 18398
rect 29038 18386 29090 18398
rect 30494 18450 30546 18462
rect 30494 18386 30546 18398
rect 32174 18450 32226 18462
rect 33282 18398 33294 18450
rect 33346 18398 33358 18450
rect 32174 18386 32226 18398
rect 2494 18338 2546 18350
rect 7646 18338 7698 18350
rect 6626 18286 6638 18338
rect 6690 18286 6702 18338
rect 2494 18274 2546 18286
rect 7646 18274 7698 18286
rect 8094 18338 8146 18350
rect 8094 18274 8146 18286
rect 10670 18338 10722 18350
rect 10670 18274 10722 18286
rect 17614 18338 17666 18350
rect 23774 18338 23826 18350
rect 29822 18338 29874 18350
rect 19282 18286 19294 18338
rect 19346 18286 19358 18338
rect 21410 18286 21422 18338
rect 21474 18286 21486 18338
rect 24546 18286 24558 18338
rect 24610 18286 24622 18338
rect 17614 18274 17666 18286
rect 23774 18274 23826 18286
rect 29822 18274 29874 18286
rect 31390 18338 31442 18350
rect 32510 18338 32562 18350
rect 31826 18286 31838 18338
rect 31890 18286 31902 18338
rect 31390 18274 31442 18286
rect 32510 18274 32562 18286
rect 18062 18226 18114 18238
rect 6066 18174 6078 18226
rect 6130 18174 6142 18226
rect 7186 18174 7198 18226
rect 7250 18223 7262 18226
rect 7634 18223 7646 18226
rect 7250 18177 7646 18223
rect 7250 18174 7262 18177
rect 7634 18174 7646 18177
rect 7698 18223 7710 18226
rect 8194 18223 8206 18226
rect 7698 18177 8206 18223
rect 7698 18174 7710 18177
rect 8194 18174 8206 18177
rect 8258 18174 8270 18226
rect 18062 18162 18114 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 30146 17838 30158 17890
rect 30210 17838 30222 17890
rect 9774 17778 9826 17790
rect 5058 17726 5070 17778
rect 5122 17726 5134 17778
rect 8082 17726 8094 17778
rect 8146 17726 8158 17778
rect 9774 17714 9826 17726
rect 19406 17778 19458 17790
rect 19406 17714 19458 17726
rect 20750 17778 20802 17790
rect 20750 17714 20802 17726
rect 25342 17778 25394 17790
rect 25342 17714 25394 17726
rect 25678 17778 25730 17790
rect 25678 17714 25730 17726
rect 27022 17778 27074 17790
rect 27022 17714 27074 17726
rect 32846 17778 32898 17790
rect 32846 17714 32898 17726
rect 7198 17666 7250 17678
rect 19182 17666 19234 17678
rect 2258 17614 2270 17666
rect 2322 17614 2334 17666
rect 7858 17614 7870 17666
rect 7922 17614 7934 17666
rect 18386 17614 18398 17666
rect 18450 17614 18462 17666
rect 7198 17602 7250 17614
rect 19182 17602 19234 17614
rect 19518 17666 19570 17678
rect 19518 17602 19570 17614
rect 19742 17666 19794 17678
rect 27246 17666 27298 17678
rect 26114 17614 26126 17666
rect 26178 17614 26190 17666
rect 19742 17602 19794 17614
rect 27246 17602 27298 17614
rect 29486 17666 29538 17678
rect 29486 17602 29538 17614
rect 29934 17666 29986 17678
rect 29934 17602 29986 17614
rect 31278 17666 31330 17678
rect 31278 17602 31330 17614
rect 31614 17666 31666 17678
rect 31614 17602 31666 17614
rect 35982 17666 36034 17678
rect 35982 17602 36034 17614
rect 6078 17554 6130 17566
rect 2930 17502 2942 17554
rect 2994 17502 3006 17554
rect 6078 17490 6130 17502
rect 6190 17554 6242 17566
rect 6190 17490 6242 17502
rect 6414 17554 6466 17566
rect 6414 17490 6466 17502
rect 6638 17554 6690 17566
rect 6638 17490 6690 17502
rect 6750 17554 6802 17566
rect 6750 17490 6802 17502
rect 6974 17554 7026 17566
rect 8430 17554 8482 17566
rect 8194 17502 8206 17554
rect 8258 17502 8270 17554
rect 6974 17490 7026 17502
rect 8430 17490 8482 17502
rect 8654 17554 8706 17566
rect 8654 17490 8706 17502
rect 8766 17554 8818 17566
rect 8766 17490 8818 17502
rect 9214 17554 9266 17566
rect 9214 17490 9266 17502
rect 9326 17554 9378 17566
rect 20302 17554 20354 17566
rect 15026 17502 15038 17554
rect 15090 17502 15102 17554
rect 9326 17490 9378 17502
rect 20302 17490 20354 17502
rect 27470 17554 27522 17566
rect 27470 17490 27522 17502
rect 27582 17554 27634 17566
rect 27582 17490 27634 17502
rect 30606 17554 30658 17566
rect 30606 17490 30658 17502
rect 30718 17554 30770 17566
rect 30718 17490 30770 17502
rect 31950 17554 32002 17566
rect 31950 17490 32002 17502
rect 5742 17442 5794 17454
rect 5742 17378 5794 17390
rect 8990 17442 9042 17454
rect 28590 17442 28642 17454
rect 28242 17390 28254 17442
rect 28306 17390 28318 17442
rect 8990 17378 9042 17390
rect 28590 17378 28642 17390
rect 30942 17442 30994 17454
rect 30942 17378 30994 17390
rect 31614 17442 31666 17454
rect 31614 17378 31666 17390
rect 36094 17442 36146 17454
rect 36094 17378 36146 17390
rect 36318 17442 36370 17454
rect 36318 17378 36370 17390
rect 37102 17442 37154 17454
rect 37102 17378 37154 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 7758 17106 7810 17118
rect 7758 17042 7810 17054
rect 8542 17106 8594 17118
rect 8542 17042 8594 17054
rect 9102 17106 9154 17118
rect 9102 17042 9154 17054
rect 11006 17106 11058 17118
rect 11006 17042 11058 17054
rect 18622 17106 18674 17118
rect 18622 17042 18674 17054
rect 19406 17106 19458 17118
rect 19406 17042 19458 17054
rect 19854 17106 19906 17118
rect 19854 17042 19906 17054
rect 21310 17106 21362 17118
rect 21310 17042 21362 17054
rect 29150 17106 29202 17118
rect 29150 17042 29202 17054
rect 30382 17106 30434 17118
rect 30382 17042 30434 17054
rect 30942 17106 30994 17118
rect 30942 17042 30994 17054
rect 31166 17106 31218 17118
rect 31166 17042 31218 17054
rect 31502 17106 31554 17118
rect 31502 17042 31554 17054
rect 33742 17106 33794 17118
rect 33742 17042 33794 17054
rect 37662 17106 37714 17118
rect 37662 17042 37714 17054
rect 6750 16994 6802 17006
rect 4050 16942 4062 16994
rect 4114 16942 4126 16994
rect 6750 16930 6802 16942
rect 6862 16994 6914 17006
rect 6862 16930 6914 16942
rect 7086 16994 7138 17006
rect 7086 16930 7138 16942
rect 7534 16994 7586 17006
rect 19742 16994 19794 17006
rect 10658 16942 10670 16994
rect 10722 16942 10734 16994
rect 18946 16942 18958 16994
rect 19010 16942 19022 16994
rect 7534 16930 7586 16942
rect 19742 16930 19794 16942
rect 20078 16994 20130 17006
rect 20078 16930 20130 16942
rect 20302 16994 20354 17006
rect 20302 16930 20354 16942
rect 20750 16994 20802 17006
rect 20750 16930 20802 16942
rect 20862 16994 20914 17006
rect 30830 16994 30882 17006
rect 22530 16942 22542 16994
rect 22594 16942 22606 16994
rect 20862 16930 20914 16942
rect 30830 16930 30882 16942
rect 33182 16994 33234 17006
rect 33182 16930 33234 16942
rect 35534 16994 35586 17006
rect 35534 16930 35586 16942
rect 36206 16994 36258 17006
rect 36206 16930 36258 16942
rect 2270 16882 2322 16894
rect 7198 16882 7250 16894
rect 1810 16830 1822 16882
rect 1874 16830 1886 16882
rect 3378 16830 3390 16882
rect 3442 16830 3454 16882
rect 2270 16818 2322 16830
rect 7198 16818 7250 16830
rect 7870 16882 7922 16894
rect 7870 16818 7922 16830
rect 20638 16882 20690 16894
rect 20638 16818 20690 16830
rect 21086 16882 21138 16894
rect 21086 16818 21138 16830
rect 21422 16882 21474 16894
rect 25454 16882 25506 16894
rect 21858 16830 21870 16882
rect 21922 16830 21934 16882
rect 21422 16818 21474 16830
rect 25454 16818 25506 16830
rect 33070 16882 33122 16894
rect 33070 16818 33122 16830
rect 33406 16882 33458 16894
rect 33406 16818 33458 16830
rect 35422 16882 35474 16894
rect 35422 16818 35474 16830
rect 35982 16882 36034 16894
rect 35982 16818 36034 16830
rect 36430 16882 36482 16894
rect 36430 16818 36482 16830
rect 36654 16882 36706 16894
rect 36654 16818 36706 16830
rect 37214 16882 37266 16894
rect 37214 16818 37266 16830
rect 35758 16770 35810 16782
rect 6178 16718 6190 16770
rect 6242 16718 6254 16770
rect 24658 16718 24670 16770
rect 24722 16718 24734 16770
rect 35758 16706 35810 16718
rect 36318 16770 36370 16782
rect 36318 16706 36370 16718
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 35982 16322 36034 16334
rect 35982 16258 36034 16270
rect 1822 16210 1874 16222
rect 1822 16146 1874 16158
rect 5742 16210 5794 16222
rect 5742 16146 5794 16158
rect 14366 16210 14418 16222
rect 14366 16146 14418 16158
rect 16158 16210 16210 16222
rect 16158 16146 16210 16158
rect 17054 16210 17106 16222
rect 17054 16146 17106 16158
rect 17950 16210 18002 16222
rect 17950 16146 18002 16158
rect 20078 16210 20130 16222
rect 20078 16146 20130 16158
rect 21646 16210 21698 16222
rect 34862 16210 34914 16222
rect 32722 16158 32734 16210
rect 32786 16158 32798 16210
rect 21646 16146 21698 16158
rect 34862 16146 34914 16158
rect 35534 16210 35586 16222
rect 37762 16158 37774 16210
rect 37826 16158 37838 16210
rect 40002 16158 40014 16210
rect 40066 16158 40078 16210
rect 35534 16146 35586 16158
rect 6078 16098 6130 16110
rect 6078 16034 6130 16046
rect 6974 16098 7026 16110
rect 6974 16034 7026 16046
rect 7198 16098 7250 16110
rect 7198 16034 7250 16046
rect 7870 16098 7922 16110
rect 7870 16034 7922 16046
rect 8206 16098 8258 16110
rect 12910 16098 12962 16110
rect 9986 16046 9998 16098
rect 10050 16046 10062 16098
rect 8206 16034 8258 16046
rect 12910 16034 12962 16046
rect 13806 16098 13858 16110
rect 13806 16034 13858 16046
rect 17390 16098 17442 16110
rect 17390 16034 17442 16046
rect 31726 16098 31778 16110
rect 36094 16098 36146 16110
rect 32050 16046 32062 16098
rect 32114 16046 32126 16098
rect 36978 16046 36990 16098
rect 37042 16046 37054 16098
rect 31726 16034 31778 16046
rect 36094 16034 36146 16046
rect 6190 15986 6242 15998
rect 6190 15922 6242 15934
rect 6414 15986 6466 15998
rect 6414 15922 6466 15934
rect 6638 15986 6690 15998
rect 6638 15922 6690 15934
rect 8094 15986 8146 15998
rect 8094 15922 8146 15934
rect 8654 15986 8706 15998
rect 14702 15986 14754 15998
rect 9762 15934 9774 15986
rect 9826 15934 9838 15986
rect 8654 15922 8706 15934
rect 14702 15922 14754 15934
rect 14814 15986 14866 15998
rect 14814 15922 14866 15934
rect 15262 15986 15314 15998
rect 15262 15922 15314 15934
rect 15374 15986 15426 15998
rect 15374 15922 15426 15934
rect 31390 15986 31442 15998
rect 31390 15922 31442 15934
rect 31502 15986 31554 15998
rect 31502 15922 31554 15934
rect 5182 15874 5234 15886
rect 5182 15810 5234 15822
rect 6750 15874 6802 15886
rect 6750 15810 6802 15822
rect 7646 15874 7698 15886
rect 7646 15810 7698 15822
rect 13470 15874 13522 15886
rect 13470 15810 13522 15822
rect 15038 15874 15090 15886
rect 15038 15810 15090 15822
rect 15598 15874 15650 15886
rect 15598 15810 15650 15822
rect 16494 15874 16546 15886
rect 31166 15874 31218 15886
rect 20626 15822 20638 15874
rect 20690 15871 20702 15874
rect 20850 15871 20862 15874
rect 20690 15825 20862 15871
rect 20690 15822 20702 15825
rect 20850 15822 20862 15825
rect 20914 15822 20926 15874
rect 16494 15810 16546 15822
rect 31166 15810 31218 15822
rect 35982 15874 36034 15886
rect 35982 15810 36034 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 6862 15538 6914 15550
rect 6862 15474 6914 15486
rect 7422 15538 7474 15550
rect 7422 15474 7474 15486
rect 7758 15538 7810 15550
rect 12798 15538 12850 15550
rect 9538 15486 9550 15538
rect 9602 15486 9614 15538
rect 12450 15486 12462 15538
rect 12514 15486 12526 15538
rect 7758 15474 7810 15486
rect 12798 15474 12850 15486
rect 13246 15538 13298 15550
rect 13246 15474 13298 15486
rect 17502 15538 17554 15550
rect 17502 15474 17554 15486
rect 19854 15538 19906 15550
rect 20638 15538 20690 15550
rect 20290 15486 20302 15538
rect 20354 15486 20366 15538
rect 19854 15474 19906 15486
rect 20638 15474 20690 15486
rect 26014 15538 26066 15550
rect 26014 15474 26066 15486
rect 29934 15538 29986 15550
rect 29934 15474 29986 15486
rect 30270 15538 30322 15550
rect 30270 15474 30322 15486
rect 31726 15538 31778 15550
rect 31726 15474 31778 15486
rect 31950 15538 32002 15550
rect 31950 15474 32002 15486
rect 39902 15538 39954 15550
rect 39902 15474 39954 15486
rect 10334 15426 10386 15438
rect 3154 15374 3166 15426
rect 3218 15374 3230 15426
rect 6178 15374 6190 15426
rect 6242 15374 6254 15426
rect 10334 15362 10386 15374
rect 10446 15426 10498 15438
rect 10446 15362 10498 15374
rect 13134 15426 13186 15438
rect 13134 15362 13186 15374
rect 19742 15426 19794 15438
rect 19742 15362 19794 15374
rect 21646 15426 21698 15438
rect 21646 15362 21698 15374
rect 21982 15426 22034 15438
rect 21982 15362 22034 15374
rect 22094 15426 22146 15438
rect 37090 15374 37102 15426
rect 37154 15374 37166 15426
rect 22094 15362 22146 15374
rect 9886 15314 9938 15326
rect 2482 15262 2494 15314
rect 2546 15262 2558 15314
rect 6290 15262 6302 15314
rect 6354 15262 6366 15314
rect 9886 15250 9938 15262
rect 10110 15314 10162 15326
rect 20974 15314 21026 15326
rect 14018 15262 14030 15314
rect 14082 15262 14094 15314
rect 10110 15250 10162 15262
rect 20974 15250 21026 15262
rect 21422 15314 21474 15326
rect 21422 15250 21474 15262
rect 22318 15314 22370 15326
rect 22318 15250 22370 15262
rect 22654 15314 22706 15326
rect 28590 15314 28642 15326
rect 26786 15262 26798 15314
rect 26850 15262 26862 15314
rect 22654 15250 22706 15262
rect 28590 15250 28642 15262
rect 30158 15314 30210 15326
rect 30158 15250 30210 15262
rect 30494 15314 30546 15326
rect 36306 15262 36318 15314
rect 36370 15262 36382 15314
rect 30494 15250 30546 15262
rect 1822 15202 1874 15214
rect 10894 15202 10946 15214
rect 19406 15202 19458 15214
rect 5282 15150 5294 15202
rect 5346 15150 5358 15202
rect 5618 15150 5630 15202
rect 5682 15150 5694 15202
rect 14690 15150 14702 15202
rect 14754 15150 14766 15202
rect 16818 15150 16830 15202
rect 16882 15150 16894 15202
rect 1822 15138 1874 15150
rect 10894 15138 10946 15150
rect 19406 15138 19458 15150
rect 21198 15202 21250 15214
rect 39230 15202 39282 15214
rect 26450 15150 26462 15202
rect 26514 15150 26526 15202
rect 32386 15150 32398 15202
rect 32450 15150 32462 15202
rect 21198 15138 21250 15150
rect 39230 15138 39282 15150
rect 13246 15090 13298 15102
rect 13246 15026 13298 15038
rect 19854 15090 19906 15102
rect 19854 15026 19906 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 19966 14754 20018 14766
rect 19966 14690 20018 14702
rect 5854 14642 5906 14654
rect 5854 14578 5906 14590
rect 6302 14642 6354 14654
rect 6302 14578 6354 14590
rect 12014 14642 12066 14654
rect 12014 14578 12066 14590
rect 14814 14642 14866 14654
rect 14814 14578 14866 14590
rect 18286 14642 18338 14654
rect 27122 14590 27134 14642
rect 27186 14590 27198 14642
rect 18286 14578 18338 14590
rect 1710 14530 1762 14542
rect 1710 14466 1762 14478
rect 2270 14530 2322 14542
rect 2270 14466 2322 14478
rect 9326 14530 9378 14542
rect 12574 14530 12626 14542
rect 10994 14478 11006 14530
rect 11058 14478 11070 14530
rect 9326 14466 9378 14478
rect 12574 14466 12626 14478
rect 14366 14530 14418 14542
rect 14366 14466 14418 14478
rect 14590 14530 14642 14542
rect 14590 14466 14642 14478
rect 15038 14530 15090 14542
rect 15038 14466 15090 14478
rect 18846 14530 18898 14542
rect 18846 14466 18898 14478
rect 19854 14530 19906 14542
rect 19854 14466 19906 14478
rect 21198 14530 21250 14542
rect 21198 14466 21250 14478
rect 21646 14530 21698 14542
rect 21646 14466 21698 14478
rect 21870 14530 21922 14542
rect 27582 14530 27634 14542
rect 26114 14478 26126 14530
rect 26178 14478 26190 14530
rect 21870 14466 21922 14478
rect 27582 14466 27634 14478
rect 28030 14530 28082 14542
rect 30146 14478 30158 14530
rect 30210 14478 30222 14530
rect 28030 14466 28082 14478
rect 12462 14418 12514 14430
rect 12462 14354 12514 14366
rect 15262 14418 15314 14430
rect 18734 14418 18786 14430
rect 16258 14366 16270 14418
rect 16322 14366 16334 14418
rect 28366 14418 28418 14430
rect 48190 14418 48242 14430
rect 15262 14354 15314 14366
rect 18734 14354 18786 14366
rect 20414 14362 20466 14374
rect 8990 14306 9042 14318
rect 8990 14242 9042 14254
rect 9438 14306 9490 14318
rect 9438 14242 9490 14254
rect 9662 14306 9714 14318
rect 9662 14242 9714 14254
rect 11230 14306 11282 14318
rect 11230 14242 11282 14254
rect 12238 14306 12290 14318
rect 12238 14242 12290 14254
rect 13918 14306 13970 14318
rect 13918 14242 13970 14254
rect 14030 14306 14082 14318
rect 14030 14242 14082 14254
rect 14254 14306 14306 14318
rect 14254 14242 14306 14254
rect 15934 14306 15986 14318
rect 15934 14242 15986 14254
rect 18510 14306 18562 14318
rect 18510 14242 18562 14254
rect 19630 14306 19682 14318
rect 19630 14242 19682 14254
rect 19966 14306 20018 14318
rect 32050 14366 32062 14418
rect 32114 14366 32126 14418
rect 28366 14354 28418 14366
rect 48190 14354 48242 14366
rect 20414 14298 20466 14310
rect 20526 14306 20578 14318
rect 19966 14242 20018 14254
rect 20526 14242 20578 14254
rect 20750 14306 20802 14318
rect 20750 14242 20802 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 25678 14306 25730 14318
rect 26686 14306 26738 14318
rect 26338 14254 26350 14306
rect 26402 14254 26414 14306
rect 25678 14242 25730 14254
rect 26686 14242 26738 14254
rect 47630 14306 47682 14318
rect 47630 14242 47682 14254
rect 47854 14306 47906 14318
rect 47854 14242 47906 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 11454 13970 11506 13982
rect 11454 13906 11506 13918
rect 27246 13970 27298 13982
rect 27246 13906 27298 13918
rect 27918 13970 27970 13982
rect 27918 13906 27970 13918
rect 28926 13970 28978 13982
rect 28926 13906 28978 13918
rect 29374 13970 29426 13982
rect 29374 13906 29426 13918
rect 9550 13858 9602 13870
rect 9550 13794 9602 13806
rect 9886 13858 9938 13870
rect 9886 13794 9938 13806
rect 10446 13858 10498 13870
rect 10446 13794 10498 13806
rect 10782 13858 10834 13870
rect 28030 13858 28082 13870
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 10782 13794 10834 13806
rect 28030 13794 28082 13806
rect 28478 13858 28530 13870
rect 28478 13794 28530 13806
rect 29822 13858 29874 13870
rect 29822 13794 29874 13806
rect 30046 13858 30098 13870
rect 30046 13794 30098 13806
rect 30270 13858 30322 13870
rect 30270 13794 30322 13806
rect 30830 13858 30882 13870
rect 30830 13794 30882 13806
rect 2270 13746 2322 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 2270 13682 2322 13694
rect 10110 13746 10162 13758
rect 10110 13682 10162 13694
rect 20862 13746 20914 13758
rect 27694 13746 27746 13758
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 20862 13682 20914 13694
rect 27694 13682 27746 13694
rect 29710 13746 29762 13758
rect 29710 13682 29762 13694
rect 30494 13746 30546 13758
rect 30494 13682 30546 13694
rect 31054 13746 31106 13758
rect 31054 13682 31106 13694
rect 31390 13746 31442 13758
rect 31390 13682 31442 13694
rect 31614 13746 31666 13758
rect 31614 13682 31666 13694
rect 9662 13634 9714 13646
rect 9662 13570 9714 13582
rect 21534 13634 21586 13646
rect 30382 13634 30434 13646
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 21534 13570 21586 13582
rect 30382 13570 30434 13582
rect 31278 13634 31330 13646
rect 31278 13570 31330 13582
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 1822 13074 1874 13086
rect 28590 13074 28642 13086
rect 34862 13074 34914 13086
rect 20290 13022 20302 13074
rect 20354 13022 20366 13074
rect 24210 13022 24222 13074
rect 24274 13022 24286 13074
rect 26338 13022 26350 13074
rect 26402 13022 26414 13074
rect 32722 13022 32734 13074
rect 32786 13022 32798 13074
rect 1822 13010 1874 13022
rect 28590 13010 28642 13022
rect 34862 13010 34914 13022
rect 11454 12962 11506 12974
rect 11454 12898 11506 12910
rect 11678 12962 11730 12974
rect 11678 12898 11730 12910
rect 12686 12962 12738 12974
rect 12686 12898 12738 12910
rect 13022 12962 13074 12974
rect 13022 12898 13074 12910
rect 13358 12962 13410 12974
rect 13358 12898 13410 12910
rect 13694 12962 13746 12974
rect 13694 12898 13746 12910
rect 13918 12962 13970 12974
rect 13918 12898 13970 12910
rect 14590 12962 14642 12974
rect 21534 12962 21586 12974
rect 27806 12962 27858 12974
rect 16706 12910 16718 12962
rect 16770 12910 16782 12962
rect 23538 12910 23550 12962
rect 23602 12910 23614 12962
rect 14590 12898 14642 12910
rect 21534 12898 21586 12910
rect 27806 12898 27858 12910
rect 29262 12962 29314 12974
rect 29262 12898 29314 12910
rect 30046 12962 30098 12974
rect 30046 12898 30098 12910
rect 30718 12962 30770 12974
rect 32050 12910 32062 12962
rect 32114 12910 32126 12962
rect 30718 12898 30770 12910
rect 11902 12850 11954 12862
rect 11902 12786 11954 12798
rect 14478 12850 14530 12862
rect 14478 12786 14530 12798
rect 27246 12850 27298 12862
rect 27246 12786 27298 12798
rect 29374 12850 29426 12862
rect 29374 12786 29426 12798
rect 30382 12850 30434 12862
rect 30382 12786 30434 12798
rect 11790 12738 11842 12750
rect 11790 12674 11842 12686
rect 12462 12738 12514 12750
rect 12462 12674 12514 12686
rect 12798 12738 12850 12750
rect 12798 12674 12850 12686
rect 13582 12738 13634 12750
rect 13582 12674 13634 12686
rect 14254 12738 14306 12750
rect 14254 12674 14306 12686
rect 26798 12738 26850 12750
rect 26798 12674 26850 12686
rect 27470 12738 27522 12750
rect 27470 12674 27522 12686
rect 27694 12738 27746 12750
rect 27694 12674 27746 12686
rect 29598 12738 29650 12750
rect 29598 12674 29650 12686
rect 29710 12738 29762 12750
rect 29710 12674 29762 12686
rect 29934 12738 29986 12750
rect 29934 12674 29986 12686
rect 30494 12738 30546 12750
rect 30494 12674 30546 12686
rect 31054 12738 31106 12750
rect 31054 12674 31106 12686
rect 31502 12738 31554 12750
rect 31502 12674 31554 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 11678 12402 11730 12414
rect 11678 12338 11730 12350
rect 11902 12402 11954 12414
rect 11902 12338 11954 12350
rect 12126 12402 12178 12414
rect 12126 12338 12178 12350
rect 14814 12402 14866 12414
rect 14814 12338 14866 12350
rect 27694 12402 27746 12414
rect 27694 12338 27746 12350
rect 12238 12290 12290 12302
rect 8194 12238 8206 12290
rect 8258 12238 8270 12290
rect 12238 12226 12290 12238
rect 13358 12290 13410 12302
rect 13358 12226 13410 12238
rect 13582 12290 13634 12302
rect 13582 12226 13634 12238
rect 18958 12290 19010 12302
rect 18958 12226 19010 12238
rect 20526 12290 20578 12302
rect 20526 12226 20578 12238
rect 27470 12290 27522 12302
rect 27470 12226 27522 12238
rect 29822 12290 29874 12302
rect 29822 12226 29874 12238
rect 14030 12178 14082 12190
rect 1810 12126 1822 12178
rect 1874 12126 1886 12178
rect 8978 12126 8990 12178
rect 9042 12126 9054 12178
rect 14030 12114 14082 12126
rect 18846 12178 18898 12190
rect 18846 12114 18898 12126
rect 19294 12178 19346 12190
rect 27694 12178 27746 12190
rect 20738 12126 20750 12178
rect 20802 12126 20814 12178
rect 19294 12114 19346 12126
rect 27694 12114 27746 12126
rect 27918 12178 27970 12190
rect 27918 12114 27970 12126
rect 28590 12178 28642 12190
rect 28590 12114 28642 12126
rect 29262 12178 29314 12190
rect 29262 12114 29314 12126
rect 29598 12178 29650 12190
rect 29598 12114 29650 12126
rect 30382 12178 30434 12190
rect 30382 12114 30434 12126
rect 2270 12066 2322 12078
rect 2270 12002 2322 12014
rect 6078 12066 6130 12078
rect 6078 12002 6130 12014
rect 9662 12066 9714 12078
rect 9662 12002 9714 12014
rect 13806 12066 13858 12078
rect 13806 12002 13858 12014
rect 19182 12066 19234 12078
rect 19182 12002 19234 12014
rect 29710 12066 29762 12078
rect 29710 12002 29762 12014
rect 31614 12066 31666 12078
rect 31614 12002 31666 12014
rect 28130 11902 28142 11954
rect 28194 11951 28206 11954
rect 28466 11951 28478 11954
rect 28194 11905 28478 11951
rect 28194 11902 28206 11905
rect 28466 11902 28478 11905
rect 28530 11902 28542 11954
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 21646 11618 21698 11630
rect 21646 11554 21698 11566
rect 1822 11506 1874 11518
rect 1822 11442 1874 11454
rect 14814 11506 14866 11518
rect 14814 11442 14866 11454
rect 16494 11506 16546 11518
rect 18050 11454 18062 11506
rect 18114 11454 18126 11506
rect 20178 11454 20190 11506
rect 20242 11454 20254 11506
rect 21970 11454 21982 11506
rect 22034 11454 22046 11506
rect 33954 11454 33966 11506
rect 34018 11454 34030 11506
rect 16494 11442 16546 11454
rect 15598 11394 15650 11406
rect 16942 11394 16994 11406
rect 20750 11394 20802 11406
rect 15810 11342 15822 11394
rect 15874 11342 15886 11394
rect 17378 11342 17390 11394
rect 17442 11342 17454 11394
rect 30930 11342 30942 11394
rect 30994 11342 31006 11394
rect 31714 11342 31726 11394
rect 31778 11342 31790 11394
rect 15598 11330 15650 11342
rect 16942 11330 16994 11342
rect 20750 11330 20802 11342
rect 15934 11282 15986 11294
rect 15934 11218 15986 11230
rect 21870 11282 21922 11294
rect 21870 11218 21922 11230
rect 34526 11170 34578 11182
rect 34526 11106 34578 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 14926 10834 14978 10846
rect 14926 10770 14978 10782
rect 16494 10834 16546 10846
rect 16494 10770 16546 10782
rect 19182 10834 19234 10846
rect 19182 10770 19234 10782
rect 20078 10834 20130 10846
rect 20078 10770 20130 10782
rect 20638 10834 20690 10846
rect 20638 10770 20690 10782
rect 20974 10834 21026 10846
rect 26226 10782 26238 10834
rect 26290 10782 26302 10834
rect 20974 10770 21026 10782
rect 2270 10722 2322 10734
rect 19406 10722 19458 10734
rect 13682 10670 13694 10722
rect 13746 10670 13758 10722
rect 2270 10658 2322 10670
rect 19406 10658 19458 10670
rect 21198 10722 21250 10734
rect 21858 10670 21870 10722
rect 21922 10670 21934 10722
rect 28466 10670 28478 10722
rect 28530 10670 28542 10722
rect 21198 10658 21250 10670
rect 19518 10610 19570 10622
rect 1810 10558 1822 10610
rect 1874 10558 1886 10610
rect 14466 10558 14478 10610
rect 14530 10558 14542 10610
rect 15362 10558 15374 10610
rect 15426 10558 15438 10610
rect 15810 10558 15822 10610
rect 15874 10558 15886 10610
rect 21634 10558 21646 10610
rect 21698 10558 21710 10610
rect 29138 10558 29150 10610
rect 29202 10558 29214 10610
rect 19518 10546 19570 10558
rect 29710 10498 29762 10510
rect 11554 10446 11566 10498
rect 11618 10446 11630 10498
rect 29710 10434 29762 10446
rect 20862 10386 20914 10398
rect 15362 10334 15374 10386
rect 15426 10334 15438 10386
rect 20862 10322 20914 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 20302 10050 20354 10062
rect 20302 9986 20354 9998
rect 22318 10050 22370 10062
rect 22318 9986 22370 9998
rect 1822 9938 1874 9950
rect 12126 9938 12178 9950
rect 9426 9886 9438 9938
rect 9490 9886 9502 9938
rect 11554 9886 11566 9938
rect 11618 9886 11630 9938
rect 1822 9874 1874 9886
rect 12126 9874 12178 9886
rect 15374 9938 15426 9950
rect 23102 9938 23154 9950
rect 32734 9938 32786 9950
rect 19954 9886 19966 9938
rect 20018 9886 20030 9938
rect 29922 9886 29934 9938
rect 29986 9886 29998 9938
rect 15374 9874 15426 9886
rect 23102 9874 23154 9886
rect 32734 9874 32786 9886
rect 14366 9826 14418 9838
rect 8754 9774 8766 9826
rect 8818 9774 8830 9826
rect 12450 9774 12462 9826
rect 12514 9774 12526 9826
rect 14130 9774 14142 9826
rect 14194 9774 14206 9826
rect 14366 9762 14418 9774
rect 15710 9826 15762 9838
rect 15710 9762 15762 9774
rect 21870 9826 21922 9838
rect 21870 9762 21922 9774
rect 22206 9826 22258 9838
rect 23550 9826 23602 9838
rect 22418 9774 22430 9826
rect 22482 9774 22494 9826
rect 22206 9762 22258 9774
rect 23550 9762 23602 9774
rect 24334 9826 24386 9838
rect 29138 9774 29150 9826
rect 29202 9774 29214 9826
rect 24334 9762 24386 9774
rect 13582 9714 13634 9726
rect 13582 9650 13634 9662
rect 24446 9714 24498 9726
rect 24446 9650 24498 9662
rect 12574 9602 12626 9614
rect 12574 9538 12626 9550
rect 14814 9602 14866 9614
rect 14814 9538 14866 9550
rect 19630 9602 19682 9614
rect 19630 9538 19682 9550
rect 20078 9602 20130 9614
rect 20078 9538 20130 9550
rect 22654 9602 22706 9614
rect 32162 9550 32174 9602
rect 32226 9550 32238 9602
rect 22654 9538 22706 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 2046 9266 2098 9278
rect 2046 9202 2098 9214
rect 11454 9266 11506 9278
rect 11454 9202 11506 9214
rect 11790 9266 11842 9278
rect 11790 9202 11842 9214
rect 12350 9266 12402 9278
rect 12350 9202 12402 9214
rect 15934 9266 15986 9278
rect 15934 9202 15986 9214
rect 18622 9266 18674 9278
rect 18622 9202 18674 9214
rect 20078 9266 20130 9278
rect 20078 9202 20130 9214
rect 20190 9154 20242 9166
rect 13346 9102 13358 9154
rect 13410 9102 13422 9154
rect 19506 9102 19518 9154
rect 19570 9102 19582 9154
rect 20190 9090 20242 9102
rect 20526 9154 20578 9166
rect 22206 9154 22258 9166
rect 20738 9102 20750 9154
rect 20802 9102 20814 9154
rect 47842 9102 47854 9154
rect 47906 9102 47918 9154
rect 20526 9090 20578 9102
rect 22206 9090 22258 9102
rect 1710 9042 1762 9054
rect 19294 9042 19346 9054
rect 12674 8990 12686 9042
rect 12738 8990 12750 9042
rect 19170 8990 19182 9042
rect 19234 8990 19246 9042
rect 1710 8978 1762 8990
rect 19294 8978 19346 8990
rect 19742 9042 19794 9054
rect 19742 8978 19794 8990
rect 20974 9042 21026 9054
rect 25902 9042 25954 9054
rect 48190 9042 48242 9054
rect 21298 8990 21310 9042
rect 21362 8990 21374 9042
rect 26226 8990 26238 9042
rect 26290 8990 26302 9042
rect 20974 8978 21026 8990
rect 25902 8978 25954 8990
rect 48190 8978 48242 8990
rect 2494 8930 2546 8942
rect 19630 8930 19682 8942
rect 15474 8878 15486 8930
rect 15538 8878 15550 8930
rect 2494 8866 2546 8878
rect 19630 8866 19682 8878
rect 20638 8930 20690 8942
rect 20638 8866 20690 8878
rect 21758 8930 21810 8942
rect 21758 8866 21810 8878
rect 26686 8930 26738 8942
rect 26686 8866 26738 8878
rect 27134 8930 27186 8942
rect 27134 8866 27186 8878
rect 47630 8930 47682 8942
rect 47630 8866 47682 8878
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 20078 8370 20130 8382
rect 23650 8318 23662 8370
rect 23714 8318 23726 8370
rect 25778 8318 25790 8370
rect 25842 8318 25854 8370
rect 20078 8306 20130 8318
rect 26350 8258 26402 8270
rect 22978 8206 22990 8258
rect 23042 8206 23054 8258
rect 26350 8194 26402 8206
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 16830 7698 16882 7710
rect 2034 7646 2046 7698
rect 2098 7646 2110 7698
rect 16830 7634 16882 7646
rect 21870 7698 21922 7710
rect 21870 7634 21922 7646
rect 19506 7534 19518 7586
rect 19570 7534 19582 7586
rect 1710 7474 1762 7486
rect 20638 7474 20690 7486
rect 20178 7422 20190 7474
rect 20242 7422 20254 7474
rect 1710 7410 1762 7422
rect 20638 7410 20690 7422
rect 21086 7474 21138 7486
rect 21086 7410 21138 7422
rect 2494 7362 2546 7374
rect 17378 7310 17390 7362
rect 17442 7310 17454 7362
rect 2494 7298 2546 7310
rect 21298 7198 21310 7250
rect 21362 7198 21374 7250
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 22654 6914 22706 6926
rect 22654 6850 22706 6862
rect 23438 6914 23490 6926
rect 23438 6850 23490 6862
rect 20414 6802 20466 6814
rect 20414 6738 20466 6750
rect 22430 6802 22482 6814
rect 22430 6738 22482 6750
rect 23662 6690 23714 6702
rect 23662 6626 23714 6638
rect 24222 6690 24274 6702
rect 24222 6626 24274 6638
rect 22766 6578 22818 6590
rect 22766 6514 22818 6526
rect 23090 6414 23102 6466
rect 23154 6414 23166 6466
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 19742 6130 19794 6142
rect 19742 6066 19794 6078
rect 20850 5966 20862 6018
rect 20914 5966 20926 6018
rect 2270 5906 2322 5918
rect 1810 5854 1822 5906
rect 1874 5854 1886 5906
rect 20178 5854 20190 5906
rect 20242 5854 20254 5906
rect 2270 5842 2322 5854
rect 22978 5742 22990 5794
rect 23042 5742 23054 5794
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 1822 5234 1874 5246
rect 1822 5170 1874 5182
rect 24110 5234 24162 5246
rect 24110 5170 24162 5182
rect 22530 5070 22542 5122
rect 22594 5070 22606 5122
rect 23090 5070 23102 5122
rect 23154 5070 23166 5122
rect 22766 5010 22818 5022
rect 22766 4946 22818 4958
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 22094 4562 22146 4574
rect 2034 4510 2046 4562
rect 2098 4510 2110 4562
rect 22094 4498 22146 4510
rect 40350 4562 40402 4574
rect 47842 4510 47854 4562
rect 47906 4510 47918 4562
rect 40350 4498 40402 4510
rect 1710 4338 1762 4350
rect 48190 4338 48242 4350
rect 7074 4286 7086 4338
rect 7138 4286 7150 4338
rect 12002 4286 12014 4338
rect 12066 4286 12078 4338
rect 13346 4286 13358 4338
rect 13410 4286 13422 4338
rect 21634 4286 21646 4338
rect 21698 4286 21710 4338
rect 27122 4286 27134 4338
rect 27186 4286 27198 4338
rect 33170 4286 33182 4338
rect 33234 4286 33246 4338
rect 41234 4286 41246 4338
rect 41298 4286 41310 4338
rect 1710 4274 1762 4286
rect 48190 4274 48242 4286
rect 2494 4226 2546 4238
rect 2494 4162 2546 4174
rect 2942 4226 2994 4238
rect 2942 4162 2994 4174
rect 46958 4226 47010 4238
rect 46958 4162 47010 4174
rect 47630 4226 47682 4238
rect 47630 4162 47682 4174
rect 5182 4114 5234 4126
rect 5182 4050 5234 4062
rect 9774 4114 9826 4126
rect 9774 4050 9826 4062
rect 14030 4114 14082 4126
rect 14030 4050 14082 4062
rect 19294 4114 19346 4126
rect 19294 4050 19346 4062
rect 28142 4114 28194 4126
rect 28142 4050 28194 4062
rect 34190 4114 34242 4126
rect 34190 4050 34242 4062
rect 42254 4114 42306 4126
rect 42254 4050 42306 4062
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 17278 3666 17330 3678
rect 2706 3614 2718 3666
rect 2770 3614 2782 3666
rect 6738 3614 6750 3666
rect 6802 3614 6814 3666
rect 17278 3602 17330 3614
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 25342 3666 25394 3678
rect 25342 3602 25394 3614
rect 40014 3666 40066 3678
rect 40014 3602 40066 3614
rect 42814 3666 42866 3678
rect 42814 3602 42866 3614
rect 43822 3666 43874 3678
rect 47842 3614 47854 3666
rect 47906 3614 47918 3666
rect 43822 3602 43874 3614
rect 20078 3554 20130 3566
rect 28478 3554 28530 3566
rect 46622 3554 46674 3566
rect 4946 3502 4958 3554
rect 5010 3502 5022 3554
rect 8306 3502 8318 3554
rect 8370 3502 8382 3554
rect 12562 3502 12574 3554
rect 12626 3502 12638 3554
rect 16034 3502 16046 3554
rect 16098 3502 16110 3554
rect 19170 3502 19182 3554
rect 19234 3502 19246 3554
rect 21298 3502 21310 3554
rect 21362 3502 21374 3554
rect 27234 3502 27246 3554
rect 27298 3502 27310 3554
rect 29026 3502 29038 3554
rect 29090 3502 29102 3554
rect 32610 3502 32622 3554
rect 32674 3502 32686 3554
rect 36194 3502 36206 3554
rect 36258 3502 36270 3554
rect 37426 3502 37438 3554
rect 37490 3502 37502 3554
rect 42018 3502 42030 3554
rect 42082 3502 42094 3554
rect 45714 3502 45726 3554
rect 45778 3502 45790 3554
rect 20078 3490 20130 3502
rect 28478 3490 28530 3502
rect 46622 3490 46674 3502
rect 1710 3442 1762 3454
rect 35534 3442 35586 3454
rect 2034 3390 2046 3442
rect 2098 3390 2110 3442
rect 10770 3390 10782 3442
rect 10834 3390 10846 3442
rect 14802 3390 14814 3442
rect 14866 3390 14878 3442
rect 33730 3390 33742 3442
rect 33794 3390 33806 3442
rect 1710 3378 1762 3390
rect 35534 3378 35586 3390
rect 35982 3442 36034 3454
rect 35982 3378 36034 3390
rect 36990 3442 37042 3454
rect 47406 3442 47458 3454
rect 37202 3390 37214 3442
rect 37266 3390 37278 3442
rect 36990 3378 37042 3390
rect 47406 3378 47458 3390
rect 30046 3330 30098 3342
rect 30046 3266 30098 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 20190 46398 20242 46450
rect 20974 46398 21026 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 26238 46062 26290 46114
rect 29486 46062 29538 46114
rect 33182 46062 33234 46114
rect 36990 46062 37042 46114
rect 40798 46062 40850 46114
rect 44606 46062 44658 46114
rect 1934 45950 1986 46002
rect 6638 45950 6690 46002
rect 7198 45950 7250 46002
rect 8094 45950 8146 46002
rect 10782 45950 10834 46002
rect 13470 45950 13522 46002
rect 14814 45950 14866 46002
rect 16382 45950 16434 46002
rect 18846 45950 18898 46002
rect 20190 45950 20242 46002
rect 22878 45950 22930 46002
rect 47630 45950 47682 46002
rect 4286 45838 4338 45890
rect 4734 45838 4786 45890
rect 5630 45838 5682 45890
rect 6190 45838 6242 45890
rect 9662 45838 9714 45890
rect 11006 45838 11058 45890
rect 12238 45838 12290 45890
rect 13694 45838 13746 45890
rect 15038 45838 15090 45890
rect 17054 45838 17106 45890
rect 17726 45838 17778 45890
rect 19294 45838 19346 45890
rect 20974 45838 21026 45890
rect 21982 45838 22034 45890
rect 23326 45838 23378 45890
rect 25230 45838 25282 45890
rect 28926 45838 28978 45890
rect 32174 45838 32226 45890
rect 35982 45838 36034 45890
rect 39790 45838 39842 45890
rect 43934 45838 43986 45890
rect 48190 45838 48242 45890
rect 8766 45726 8818 45778
rect 4958 45614 5010 45666
rect 8430 45614 8482 45666
rect 9998 45614 10050 45666
rect 11342 45614 11394 45666
rect 12574 45614 12626 45666
rect 14030 45614 14082 45666
rect 15374 45614 15426 45666
rect 17278 45614 17330 45666
rect 18062 45614 18114 45666
rect 19070 45614 19122 45666
rect 20750 45614 20802 45666
rect 21758 45614 21810 45666
rect 23102 45614 23154 45666
rect 47854 45614 47906 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 9662 45278 9714 45330
rect 11678 45278 11730 45330
rect 12798 45278 12850 45330
rect 17614 45278 17666 45330
rect 21534 45278 21586 45330
rect 28142 45278 28194 45330
rect 31838 45278 31890 45330
rect 36990 45278 37042 45330
rect 41918 45278 41970 45330
rect 44830 45278 44882 45330
rect 7534 45166 7586 45218
rect 7870 45166 7922 45218
rect 8654 45166 8706 45218
rect 25902 45166 25954 45218
rect 3950 45054 4002 45106
rect 7198 45054 7250 45106
rect 8430 45054 8482 45106
rect 12014 45054 12066 45106
rect 25566 45054 25618 45106
rect 27134 45054 27186 45106
rect 31614 45054 31666 45106
rect 35198 45054 35250 45106
rect 35982 45054 36034 45106
rect 41022 45054 41074 45106
rect 43822 45054 43874 45106
rect 4846 44942 4898 44994
rect 30158 44942 30210 44994
rect 33294 44942 33346 44994
rect 1934 44830 1986 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 25454 44494 25506 44546
rect 28478 44494 28530 44546
rect 30830 44494 30882 44546
rect 37998 44494 38050 44546
rect 40910 44494 40962 44546
rect 45838 44494 45890 44546
rect 1934 44382 1986 44434
rect 8878 44382 8930 44434
rect 15262 44382 15314 44434
rect 16382 44382 16434 44434
rect 27470 44382 27522 44434
rect 27918 44382 27970 44434
rect 4846 44270 4898 44322
rect 5966 44270 6018 44322
rect 14702 44270 14754 44322
rect 19182 44270 19234 44322
rect 24446 44270 24498 44322
rect 28254 44270 28306 44322
rect 29374 44270 29426 44322
rect 29934 44270 29986 44322
rect 35422 44270 35474 44322
rect 36990 44270 37042 44322
rect 39902 44270 39954 44322
rect 44830 44270 44882 44322
rect 4062 44158 4114 44210
rect 6750 44158 6802 44210
rect 11342 44158 11394 44210
rect 18510 44158 18562 44210
rect 22430 44158 22482 44210
rect 22766 44158 22818 44210
rect 23774 44158 23826 44210
rect 24110 44158 24162 44210
rect 29150 44158 29202 44210
rect 32734 44158 32786 44210
rect 33070 44158 33122 44210
rect 33406 44158 33458 44210
rect 33742 44158 33794 44210
rect 34078 44158 34130 44210
rect 34414 44158 34466 44210
rect 35646 44158 35698 44210
rect 42814 44158 42866 44210
rect 43150 44158 43202 44210
rect 43486 44158 43538 44210
rect 43822 44158 43874 44210
rect 9326 44046 9378 44098
rect 11678 44046 11730 44098
rect 14814 44046 14866 44098
rect 15150 44046 15202 44098
rect 19742 44046 19794 44098
rect 21534 44046 21586 44098
rect 21870 44046 21922 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 5294 43710 5346 43762
rect 29934 43710 29986 43762
rect 6750 43598 6802 43650
rect 7422 43598 7474 43650
rect 8094 43598 8146 43650
rect 10558 43598 10610 43650
rect 17950 43598 18002 43650
rect 20974 43598 21026 43650
rect 31614 43598 31666 43650
rect 33406 43598 33458 43650
rect 45278 43598 45330 43650
rect 4286 43486 4338 43538
rect 4734 43486 4786 43538
rect 6974 43486 7026 43538
rect 7870 43486 7922 43538
rect 8206 43486 8258 43538
rect 10446 43486 10498 43538
rect 11342 43486 11394 43538
rect 18062 43486 18114 43538
rect 21310 43486 21362 43538
rect 25342 43486 25394 43538
rect 29598 43486 29650 43538
rect 30158 43486 30210 43538
rect 31278 43486 31330 43538
rect 33182 43486 33234 43538
rect 44942 43486 44994 43538
rect 45614 43486 45666 43538
rect 5630 43374 5682 43426
rect 12126 43374 12178 43426
rect 14254 43374 14306 43426
rect 14814 43374 14866 43426
rect 18510 43374 18562 43426
rect 19182 43374 19234 43426
rect 20414 43374 20466 43426
rect 22094 43374 22146 43426
rect 24222 43374 24274 43426
rect 26014 43374 26066 43426
rect 28142 43374 28194 43426
rect 28702 43374 28754 43426
rect 29038 43374 29090 43426
rect 44606 43374 44658 43426
rect 46622 43374 46674 43426
rect 1934 43262 1986 43314
rect 7534 43262 7586 43314
rect 10558 43262 10610 43314
rect 17950 43262 18002 43314
rect 19406 43262 19458 43314
rect 19742 43262 19794 43314
rect 20638 43262 20690 43314
rect 29262 43262 29314 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 23998 42926 24050 42978
rect 24334 42926 24386 42978
rect 41582 42926 41634 42978
rect 41918 42926 41970 42978
rect 47070 42926 47122 42978
rect 2046 42814 2098 42866
rect 12686 42814 12738 42866
rect 15038 42814 15090 42866
rect 18398 42814 18450 42866
rect 21422 42814 21474 42866
rect 22542 42814 22594 42866
rect 24782 42814 24834 42866
rect 4286 42702 4338 42754
rect 4734 42702 4786 42754
rect 8766 42702 8818 42754
rect 9886 42702 9938 42754
rect 17838 42702 17890 42754
rect 18174 42702 18226 42754
rect 22094 42702 22146 42754
rect 22318 42702 22370 42754
rect 22878 42702 22930 42754
rect 23774 42702 23826 42754
rect 28478 42702 28530 42754
rect 40910 42702 40962 42754
rect 45614 42702 45666 42754
rect 7758 42590 7810 42642
rect 8094 42590 8146 42642
rect 10558 42590 10610 42642
rect 13582 42590 13634 42642
rect 17166 42590 17218 42642
rect 18622 42590 18674 42642
rect 18846 42590 18898 42642
rect 21758 42590 21810 42642
rect 21870 42590 21922 42642
rect 22766 42590 22818 42642
rect 39790 42590 39842 42642
rect 40798 42590 40850 42642
rect 4958 42478 5010 42530
rect 8430 42478 8482 42530
rect 8654 42478 8706 42530
rect 9326 42478 9378 42530
rect 19406 42478 19458 42530
rect 19966 42478 20018 42530
rect 23438 42478 23490 42530
rect 29262 42478 29314 42530
rect 40238 42478 40290 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 10558 42142 10610 42194
rect 11790 42142 11842 42194
rect 17726 42142 17778 42194
rect 22318 42142 22370 42194
rect 7870 42030 7922 42082
rect 8430 42030 8482 42082
rect 8878 42030 8930 42082
rect 9886 42030 9938 42082
rect 9998 42030 10050 42082
rect 10222 42030 10274 42082
rect 18174 42030 18226 42082
rect 18398 42030 18450 42082
rect 18510 42030 18562 42082
rect 22206 42030 22258 42082
rect 3838 41918 3890 41970
rect 7086 41918 7138 41970
rect 7310 41918 7362 41970
rect 7646 41918 7698 41970
rect 7982 41918 8034 41970
rect 8206 41918 8258 41970
rect 8654 41918 8706 41970
rect 8990 41918 9042 41970
rect 10334 41918 10386 41970
rect 10782 41918 10834 41970
rect 10894 41918 10946 41970
rect 11342 41918 11394 41970
rect 11678 41918 11730 41970
rect 11902 41918 11954 41970
rect 16942 41918 16994 41970
rect 17390 41918 17442 41970
rect 17726 41918 17778 41970
rect 18062 41918 18114 41970
rect 22542 41918 22594 41970
rect 23214 41918 23266 41970
rect 23438 41918 23490 41970
rect 23550 41918 23602 41970
rect 23886 41918 23938 41970
rect 27918 41918 27970 41970
rect 4510 41806 4562 41858
rect 6638 41806 6690 41858
rect 7422 41806 7474 41858
rect 22878 41806 22930 41858
rect 28590 41806 28642 41858
rect 30718 41806 30770 41858
rect 31166 41806 31218 41858
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 11902 41358 11954 41410
rect 12462 41358 12514 41410
rect 18622 41358 18674 41410
rect 23214 41358 23266 41410
rect 4846 41246 4898 41298
rect 9214 41246 9266 41298
rect 23774 41246 23826 41298
rect 28030 41246 28082 41298
rect 2046 41134 2098 41186
rect 8318 41134 8370 41186
rect 12014 41134 12066 41186
rect 12574 41134 12626 41186
rect 17838 41134 17890 41186
rect 20302 41134 20354 41186
rect 22878 41134 22930 41186
rect 27582 41134 27634 41186
rect 28254 41134 28306 41186
rect 2718 41022 2770 41074
rect 8094 41022 8146 41074
rect 11566 41022 11618 41074
rect 11902 41022 11954 41074
rect 18174 41022 18226 41074
rect 18734 41022 18786 41074
rect 20078 41022 20130 41074
rect 22542 41022 22594 41074
rect 23102 41022 23154 41074
rect 27806 41022 27858 41074
rect 47630 41022 47682 41074
rect 48190 41022 48242 41074
rect 5742 40910 5794 40962
rect 6862 40910 6914 40962
rect 12462 40910 12514 40962
rect 13694 40910 13746 40962
rect 17726 40910 17778 40962
rect 18062 40910 18114 40962
rect 18622 40910 18674 40962
rect 19294 40910 19346 40962
rect 22318 40910 22370 40962
rect 22654 40910 22706 40962
rect 23214 40910 23266 40962
rect 28590 40910 28642 40962
rect 47854 40910 47906 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 8990 40574 9042 40626
rect 13022 40574 13074 40626
rect 13582 40574 13634 40626
rect 13806 40574 13858 40626
rect 14366 40574 14418 40626
rect 20414 40574 20466 40626
rect 26574 40574 26626 40626
rect 27806 40574 27858 40626
rect 28142 40574 28194 40626
rect 28366 40574 28418 40626
rect 29150 40574 29202 40626
rect 6750 40462 6802 40514
rect 7086 40462 7138 40514
rect 8430 40462 8482 40514
rect 8542 40462 8594 40514
rect 27022 40462 27074 40514
rect 27582 40462 27634 40514
rect 4286 40350 4338 40402
rect 8206 40350 8258 40402
rect 13358 40350 13410 40402
rect 13918 40350 13970 40402
rect 20638 40350 20690 40402
rect 26910 40350 26962 40402
rect 27246 40350 27298 40402
rect 27470 40350 27522 40402
rect 28030 40350 28082 40402
rect 28814 40350 28866 40402
rect 32510 40238 32562 40290
rect 1934 40126 1986 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 15038 39678 15090 39730
rect 15374 39678 15426 39730
rect 15710 39678 15762 39730
rect 16830 39678 16882 39730
rect 26126 39678 26178 39730
rect 28142 39678 28194 39730
rect 30158 39678 30210 39730
rect 32286 39678 32338 39730
rect 35534 39678 35586 39730
rect 7086 39566 7138 39618
rect 7310 39566 7362 39618
rect 14590 39566 14642 39618
rect 23326 39566 23378 39618
rect 27246 39566 27298 39618
rect 27582 39566 27634 39618
rect 27918 39566 27970 39618
rect 28254 39566 28306 39618
rect 28478 39566 28530 39618
rect 29486 39566 29538 39618
rect 32734 39566 32786 39618
rect 35982 39566 36034 39618
rect 39566 39566 39618 39618
rect 6750 39454 6802 39506
rect 14702 39454 14754 39506
rect 21982 39454 22034 39506
rect 22318 39454 22370 39506
rect 23774 39454 23826 39506
rect 23998 39454 24050 39506
rect 26462 39454 26514 39506
rect 26574 39454 26626 39506
rect 33406 39454 33458 39506
rect 6974 39342 7026 39394
rect 14142 39342 14194 39394
rect 14254 39342 14306 39394
rect 14814 39342 14866 39394
rect 16270 39342 16322 39394
rect 17390 39342 17442 39394
rect 17838 39342 17890 39394
rect 21310 39342 21362 39394
rect 21646 39342 21698 39394
rect 23662 39342 23714 39394
rect 26798 39342 26850 39394
rect 27358 39342 27410 39394
rect 39790 39342 39842 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 10222 39006 10274 39058
rect 12014 39006 12066 39058
rect 12574 39006 12626 39058
rect 13918 39006 13970 39058
rect 14478 39006 14530 39058
rect 16830 39006 16882 39058
rect 25342 39006 25394 39058
rect 27582 39006 27634 39058
rect 28366 39006 28418 39058
rect 28702 39006 28754 39058
rect 30382 39006 30434 39058
rect 32510 39006 32562 39058
rect 33966 39006 34018 39058
rect 35646 39006 35698 39058
rect 7310 38894 7362 38946
rect 14702 38894 14754 38946
rect 16718 38894 16770 38946
rect 18622 38894 18674 38946
rect 18846 38894 18898 38946
rect 23886 38894 23938 38946
rect 26910 38894 26962 38946
rect 27022 38894 27074 38946
rect 27246 38894 27298 38946
rect 27470 38894 27522 38946
rect 30942 38894 30994 38946
rect 31502 38894 31554 38946
rect 32062 38894 32114 38946
rect 34526 38894 34578 38946
rect 34974 38894 35026 38946
rect 36094 38894 36146 38946
rect 4286 38782 4338 38834
rect 8094 38782 8146 38834
rect 9886 38782 9938 38834
rect 10558 38782 10610 38834
rect 12126 38782 12178 38834
rect 12462 38782 12514 38834
rect 12798 38782 12850 38834
rect 15262 38782 15314 38834
rect 16046 38782 16098 38834
rect 16494 38782 16546 38834
rect 17502 38782 17554 38834
rect 18510 38782 18562 38834
rect 24670 38782 24722 38834
rect 27694 38782 27746 38834
rect 27918 38782 27970 38834
rect 4846 38670 4898 38722
rect 5182 38670 5234 38722
rect 8542 38670 8594 38722
rect 11454 38670 11506 38722
rect 11902 38670 11954 38722
rect 13582 38670 13634 38722
rect 17838 38670 17890 38722
rect 19182 38670 19234 38722
rect 21758 38670 21810 38722
rect 26574 38670 26626 38722
rect 30718 38670 30770 38722
rect 33294 38670 33346 38722
rect 34302 38670 34354 38722
rect 36654 38670 36706 38722
rect 1934 38558 1986 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 23326 38222 23378 38274
rect 40126 38222 40178 38274
rect 2830 38110 2882 38162
rect 3390 38110 3442 38162
rect 11118 38110 11170 38162
rect 12462 38110 12514 38162
rect 13694 38110 13746 38162
rect 16606 38110 16658 38162
rect 3278 37998 3330 38050
rect 3614 37998 3666 38050
rect 3726 37998 3778 38050
rect 3838 37998 3890 38050
rect 5182 37998 5234 38050
rect 9998 37998 10050 38050
rect 10446 37998 10498 38050
rect 18734 37998 18786 38050
rect 22430 37998 22482 38050
rect 22766 37998 22818 38050
rect 23214 37998 23266 38050
rect 29374 37998 29426 38050
rect 39006 37998 39058 38050
rect 39790 37998 39842 38050
rect 4510 37886 4562 37938
rect 4846 37886 4898 37938
rect 8094 37886 8146 37938
rect 39118 37886 39170 37938
rect 40686 37886 40738 37938
rect 2942 37774 2994 37826
rect 4398 37774 4450 37826
rect 4958 37774 5010 37826
rect 7758 37774 7810 37826
rect 10222 37774 10274 37826
rect 10334 37774 10386 37826
rect 10558 37774 10610 37826
rect 20302 37774 20354 37826
rect 22094 37774 22146 37826
rect 22542 37774 22594 37826
rect 23326 37774 23378 37826
rect 29150 37774 29202 37826
rect 41134 37774 41186 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 7646 37438 7698 37490
rect 9438 37438 9490 37490
rect 11902 37438 11954 37490
rect 13806 37438 13858 37490
rect 18622 37438 18674 37490
rect 19630 37438 19682 37490
rect 28814 37438 28866 37490
rect 29374 37438 29426 37490
rect 32510 37438 32562 37490
rect 34302 37438 34354 37490
rect 9550 37326 9602 37378
rect 11454 37326 11506 37378
rect 12462 37326 12514 37378
rect 14254 37326 14306 37378
rect 16158 37326 16210 37378
rect 17614 37326 17666 37378
rect 18062 37326 18114 37378
rect 27918 37326 27970 37378
rect 28142 37326 28194 37378
rect 33294 37326 33346 37378
rect 33742 37326 33794 37378
rect 34862 37326 34914 37378
rect 2382 37214 2434 37266
rect 5630 37214 5682 37266
rect 7982 37214 8034 37266
rect 9886 37214 9938 37266
rect 10670 37214 10722 37266
rect 10894 37214 10946 37266
rect 12686 37214 12738 37266
rect 14814 37214 14866 37266
rect 15374 37214 15426 37266
rect 15822 37214 15874 37266
rect 28478 37214 28530 37266
rect 29934 37214 29986 37266
rect 3054 37102 3106 37154
rect 5182 37102 5234 37154
rect 13246 37102 13298 37154
rect 14478 37102 14530 37154
rect 16830 37102 16882 37154
rect 19070 37102 19122 37154
rect 20078 37102 20130 37154
rect 20526 37102 20578 37154
rect 27246 37102 27298 37154
rect 33966 37102 34018 37154
rect 35422 37102 35474 37154
rect 18286 36990 18338 37042
rect 19294 36990 19346 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 4958 36654 5010 36706
rect 12014 36654 12066 36706
rect 1934 36542 1986 36594
rect 5742 36542 5794 36594
rect 11118 36542 11170 36594
rect 12238 36542 12290 36594
rect 13582 36542 13634 36594
rect 15598 36542 15650 36594
rect 19294 36542 19346 36594
rect 20302 36542 20354 36594
rect 20862 36542 20914 36594
rect 21422 36542 21474 36594
rect 32622 36542 32674 36594
rect 4286 36430 4338 36482
rect 5630 36430 5682 36482
rect 5854 36430 5906 36482
rect 6078 36430 6130 36482
rect 6414 36430 6466 36482
rect 8878 36430 8930 36482
rect 9550 36430 9602 36482
rect 9774 36430 9826 36482
rect 9998 36430 10050 36482
rect 11566 36430 11618 36482
rect 12462 36430 12514 36482
rect 13470 36430 13522 36482
rect 13694 36430 13746 36482
rect 13918 36430 13970 36482
rect 14030 36430 14082 36482
rect 15150 36430 15202 36482
rect 16606 36430 16658 36482
rect 17166 36430 17218 36482
rect 17390 36430 17442 36482
rect 18398 36430 18450 36482
rect 30046 36430 30098 36482
rect 41022 36430 41074 36482
rect 5070 36318 5122 36370
rect 8206 36318 8258 36370
rect 8430 36318 8482 36370
rect 10222 36318 10274 36370
rect 11790 36318 11842 36370
rect 16158 36318 16210 36370
rect 17950 36318 18002 36370
rect 22206 36318 22258 36370
rect 22318 36318 22370 36370
rect 47630 36318 47682 36370
rect 48190 36318 48242 36370
rect 6862 36206 6914 36258
rect 8654 36206 8706 36258
rect 9886 36206 9938 36258
rect 10670 36206 10722 36258
rect 12014 36206 12066 36258
rect 12910 36206 12962 36258
rect 14702 36206 14754 36258
rect 15934 36206 15986 36258
rect 18846 36206 18898 36258
rect 19854 36206 19906 36258
rect 21534 36206 21586 36258
rect 22542 36206 22594 36258
rect 22878 36206 22930 36258
rect 28590 36206 28642 36258
rect 41246 36206 41298 36258
rect 47854 36206 47906 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4622 35870 4674 35922
rect 9550 35870 9602 35922
rect 14814 35870 14866 35922
rect 15710 35870 15762 35922
rect 16046 35870 16098 35922
rect 16382 35870 16434 35922
rect 19182 35870 19234 35922
rect 24558 35870 24610 35922
rect 18622 35758 18674 35810
rect 19294 35758 19346 35810
rect 19742 35758 19794 35810
rect 32174 35758 32226 35810
rect 32398 35758 32450 35810
rect 4286 35646 4338 35698
rect 4958 35646 5010 35698
rect 9886 35646 9938 35698
rect 12350 35646 12402 35698
rect 14030 35646 14082 35698
rect 14366 35646 14418 35698
rect 18286 35646 18338 35698
rect 24110 35646 24162 35698
rect 33070 35646 33122 35698
rect 36430 35646 36482 35698
rect 10446 35534 10498 35586
rect 12574 35534 12626 35586
rect 15262 35534 15314 35586
rect 17502 35534 17554 35586
rect 18062 35534 18114 35586
rect 18846 35534 18898 35586
rect 19070 35534 19122 35586
rect 21198 35534 21250 35586
rect 23326 35534 23378 35586
rect 29822 35534 29874 35586
rect 31838 35534 31890 35586
rect 32510 35534 32562 35586
rect 33854 35534 33906 35586
rect 35982 35534 36034 35586
rect 37214 35534 37266 35586
rect 39342 35534 39394 35586
rect 1934 35422 1986 35474
rect 12014 35422 12066 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 4734 35086 4786 35138
rect 7310 35086 7362 35138
rect 24894 35086 24946 35138
rect 30606 35086 30658 35138
rect 34750 35086 34802 35138
rect 41246 35086 41298 35138
rect 41582 35086 41634 35138
rect 8318 34974 8370 35026
rect 13694 34974 13746 35026
rect 30270 34974 30322 35026
rect 32734 34974 32786 35026
rect 36094 34974 36146 35026
rect 2830 34862 2882 34914
rect 3278 34862 3330 34914
rect 3614 34862 3666 34914
rect 3838 34862 3890 34914
rect 4062 34862 4114 34914
rect 8990 34862 9042 34914
rect 9774 34862 9826 34914
rect 12238 34862 12290 34914
rect 18734 34862 18786 34914
rect 22430 34862 22482 34914
rect 22878 34862 22930 34914
rect 24334 34862 24386 34914
rect 24558 34862 24610 34914
rect 30046 34862 30098 34914
rect 35086 34862 35138 34914
rect 40462 34862 40514 34914
rect 2942 34750 2994 34802
rect 4398 34750 4450 34802
rect 5630 34750 5682 34802
rect 5966 34750 6018 34802
rect 7310 34750 7362 34802
rect 7422 34750 7474 34802
rect 9438 34750 9490 34802
rect 9662 34750 9714 34802
rect 12574 34750 12626 34802
rect 29150 34750 29202 34802
rect 29710 34750 29762 34802
rect 40686 34750 40738 34802
rect 42142 34750 42194 34802
rect 2382 34638 2434 34690
rect 2718 34638 2770 34690
rect 3614 34638 3666 34690
rect 4622 34638 4674 34690
rect 7870 34638 7922 34690
rect 8766 34638 8818 34690
rect 12462 34638 12514 34690
rect 12686 34638 12738 34690
rect 12798 34638 12850 34690
rect 19182 34638 19234 34690
rect 22878 34638 22930 34690
rect 29262 34638 29314 34690
rect 34862 34638 34914 34690
rect 40126 34638 40178 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2046 34302 2098 34354
rect 13134 34302 13186 34354
rect 13470 34302 13522 34354
rect 18510 34302 18562 34354
rect 25342 34302 25394 34354
rect 35534 34302 35586 34354
rect 3838 34190 3890 34242
rect 4062 34190 4114 34242
rect 12238 34190 12290 34242
rect 12350 34190 12402 34242
rect 14030 34190 14082 34242
rect 19294 34190 19346 34242
rect 19518 34190 19570 34242
rect 26126 34190 26178 34242
rect 26462 34190 26514 34242
rect 1710 34078 1762 34130
rect 12014 34078 12066 34130
rect 12462 34078 12514 34130
rect 13918 34078 13970 34130
rect 14254 34078 14306 34130
rect 18622 34078 18674 34130
rect 19070 34078 19122 34130
rect 24446 34078 24498 34130
rect 30382 34078 30434 34130
rect 35198 34078 35250 34130
rect 35534 34078 35586 34130
rect 35870 34078 35922 34130
rect 2494 33966 2546 34018
rect 3390 33966 3442 34018
rect 3726 33966 3778 34018
rect 4510 33966 4562 34018
rect 4958 33966 5010 34018
rect 18846 33966 18898 34018
rect 19966 33966 20018 34018
rect 21646 33966 21698 34018
rect 23774 33966 23826 34018
rect 26910 33966 26962 34018
rect 27470 33966 27522 34018
rect 29598 33966 29650 34018
rect 30942 33966 30994 34018
rect 4286 33854 4338 33906
rect 4622 33854 4674 33906
rect 4958 33854 5010 33906
rect 11566 33854 11618 33906
rect 30606 33854 30658 33906
rect 30942 33854 30994 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 23102 33518 23154 33570
rect 34190 33518 34242 33570
rect 34526 33518 34578 33570
rect 34974 33518 35026 33570
rect 17726 33406 17778 33458
rect 27022 33406 27074 33458
rect 28590 33406 28642 33458
rect 29262 33406 29314 33458
rect 34526 33406 34578 33458
rect 35534 33406 35586 33458
rect 38894 33406 38946 33458
rect 41022 33406 41074 33458
rect 9550 33294 9602 33346
rect 17838 33294 17890 33346
rect 18510 33294 18562 33346
rect 27694 33294 27746 33346
rect 29038 33294 29090 33346
rect 29374 33294 29426 33346
rect 30158 33294 30210 33346
rect 35310 33294 35362 33346
rect 35870 33294 35922 33346
rect 38110 33294 38162 33346
rect 9774 33182 9826 33234
rect 9886 33182 9938 33234
rect 17054 33182 17106 33234
rect 17390 33182 17442 33234
rect 22990 33182 23042 33234
rect 27358 33182 27410 33234
rect 27470 33182 27522 33234
rect 27918 33182 27970 33234
rect 28030 33182 28082 33234
rect 28254 33182 28306 33234
rect 29710 33182 29762 33234
rect 30382 33182 30434 33234
rect 10446 33070 10498 33122
rect 12910 33070 12962 33122
rect 17614 33070 17666 33122
rect 17950 33070 18002 33122
rect 22654 33070 22706 33122
rect 34862 33126 34914 33178
rect 35758 33182 35810 33234
rect 34974 33070 35026 33122
rect 37774 33070 37826 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 12014 32734 12066 32786
rect 13246 32734 13298 32786
rect 19518 32734 19570 32786
rect 26574 32734 26626 32786
rect 28366 32734 28418 32786
rect 29374 32734 29426 32786
rect 35086 32734 35138 32786
rect 10670 32622 10722 32674
rect 18174 32622 18226 32674
rect 18286 32622 18338 32674
rect 27022 32622 27074 32674
rect 27470 32622 27522 32674
rect 27582 32622 27634 32674
rect 29150 32622 29202 32674
rect 34862 32622 34914 32674
rect 35422 32622 35474 32674
rect 35646 32622 35698 32674
rect 4286 32510 4338 32562
rect 11006 32510 11058 32562
rect 12350 32510 12402 32562
rect 12910 32510 12962 32562
rect 13806 32510 13858 32562
rect 14366 32510 14418 32562
rect 18062 32510 18114 32562
rect 27134 32510 27186 32562
rect 27806 32510 27858 32562
rect 28030 32510 28082 32562
rect 28366 32510 28418 32562
rect 28702 32510 28754 32562
rect 29038 32510 29090 32562
rect 34750 32510 34802 32562
rect 35310 32510 35362 32562
rect 35870 32510 35922 32562
rect 36094 32510 36146 32562
rect 36430 32510 36482 32562
rect 37438 32510 37490 32562
rect 5070 32398 5122 32450
rect 12574 32398 12626 32450
rect 20302 32398 20354 32450
rect 29710 32398 29762 32450
rect 34414 32398 34466 32450
rect 36318 32398 36370 32450
rect 36878 32398 36930 32450
rect 38222 32398 38274 32450
rect 40350 32398 40402 32450
rect 1934 32286 1986 32338
rect 17614 32286 17666 32338
rect 27022 32286 27074 32338
rect 29486 32286 29538 32338
rect 29822 32286 29874 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 12574 31950 12626 32002
rect 1934 31838 1986 31890
rect 9102 31838 9154 31890
rect 9886 31838 9938 31890
rect 10110 31838 10162 31890
rect 10782 31838 10834 31890
rect 14926 31838 14978 31890
rect 19406 31838 19458 31890
rect 30830 31838 30882 31890
rect 4846 31726 4898 31778
rect 5742 31726 5794 31778
rect 8878 31726 8930 31778
rect 9326 31726 9378 31778
rect 10334 31726 10386 31778
rect 12126 31726 12178 31778
rect 19742 31726 19794 31778
rect 19966 31726 20018 31778
rect 31166 31726 31218 31778
rect 4062 31614 4114 31666
rect 9662 31614 9714 31666
rect 11902 31614 11954 31666
rect 12014 31614 12066 31666
rect 12686 31614 12738 31666
rect 27246 31614 27298 31666
rect 34414 31614 34466 31666
rect 5854 31502 5906 31554
rect 8318 31502 8370 31554
rect 8542 31502 8594 31554
rect 9774 31502 9826 31554
rect 11454 31502 11506 31554
rect 13582 31502 13634 31554
rect 19070 31502 19122 31554
rect 19406 31502 19458 31554
rect 19518 31502 19570 31554
rect 20526 31502 20578 31554
rect 27582 31502 27634 31554
rect 37102 31502 37154 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 7982 31166 8034 31218
rect 9438 31166 9490 31218
rect 10894 31166 10946 31218
rect 14590 31166 14642 31218
rect 18958 31166 19010 31218
rect 19070 31166 19122 31218
rect 19182 31166 19234 31218
rect 19966 31166 20018 31218
rect 22766 31166 22818 31218
rect 23214 31166 23266 31218
rect 24446 31166 24498 31218
rect 28030 31166 28082 31218
rect 33742 31166 33794 31218
rect 34190 31166 34242 31218
rect 35870 31166 35922 31218
rect 36206 31166 36258 31218
rect 36990 31166 37042 31218
rect 37998 31166 38050 31218
rect 41246 31166 41298 31218
rect 41694 31166 41746 31218
rect 43486 31166 43538 31218
rect 6078 31054 6130 31106
rect 8094 31054 8146 31106
rect 13806 31054 13858 31106
rect 14478 31054 14530 31106
rect 15262 31054 15314 31106
rect 15374 31054 15426 31106
rect 18174 31054 18226 31106
rect 20302 31054 20354 31106
rect 22318 31054 22370 31106
rect 27246 31054 27298 31106
rect 27358 31054 27410 31106
rect 27582 31054 27634 31106
rect 28366 31054 28418 31106
rect 28814 31054 28866 31106
rect 28926 31054 28978 31106
rect 34078 31054 34130 31106
rect 34862 31054 34914 31106
rect 36430 31054 36482 31106
rect 36878 31054 36930 31106
rect 42590 31054 42642 31106
rect 47854 31054 47906 31106
rect 6750 30942 6802 30994
rect 7310 30942 7362 30994
rect 7758 30942 7810 30994
rect 8766 30942 8818 30994
rect 9102 30942 9154 30994
rect 9550 30942 9602 30994
rect 9774 30942 9826 30994
rect 9998 30942 10050 30994
rect 10222 30942 10274 30994
rect 10558 30942 10610 30994
rect 13582 30942 13634 30994
rect 14030 30942 14082 30994
rect 15598 30942 15650 30994
rect 18398 30942 18450 30994
rect 19294 30942 19346 30994
rect 19518 30942 19570 30994
rect 20638 30942 20690 30994
rect 20750 30942 20802 30994
rect 21534 30942 21586 30994
rect 21758 30942 21810 30994
rect 27694 30942 27746 30994
rect 28142 30942 28194 30994
rect 28590 30942 28642 30994
rect 34750 30942 34802 30994
rect 36542 30942 36594 30994
rect 42366 30942 42418 30994
rect 43150 30942 43202 30994
rect 48190 30942 48242 30994
rect 3950 30830 4002 30882
rect 7646 30830 7698 30882
rect 8318 30830 8370 30882
rect 8542 30830 8594 30882
rect 11454 30830 11506 30882
rect 13246 30830 13298 30882
rect 14254 30830 14306 30882
rect 16046 30830 16098 30882
rect 17838 30830 17890 30882
rect 29374 30830 29426 30882
rect 37550 30830 37602 30882
rect 47630 30830 47682 30882
rect 10670 30718 10722 30770
rect 11454 30718 11506 30770
rect 14814 30718 14866 30770
rect 34190 30718 34242 30770
rect 35534 30718 35586 30770
rect 36990 30718 37042 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 25230 30382 25282 30434
rect 1934 30270 1986 30322
rect 18510 30270 18562 30322
rect 19742 30270 19794 30322
rect 20638 30270 20690 30322
rect 21646 30270 21698 30322
rect 33966 30270 34018 30322
rect 34414 30270 34466 30322
rect 41806 30270 41858 30322
rect 3950 30158 4002 30210
rect 9102 30158 9154 30210
rect 9774 30158 9826 30210
rect 14254 30158 14306 30210
rect 14702 30158 14754 30210
rect 15598 30158 15650 30210
rect 16718 30158 16770 30210
rect 24558 30158 24610 30210
rect 25006 30158 25058 30210
rect 25566 30158 25618 30210
rect 26014 30158 26066 30210
rect 30158 30158 30210 30210
rect 30382 30158 30434 30210
rect 31166 30158 31218 30210
rect 31838 30158 31890 30210
rect 35982 30158 36034 30210
rect 38894 30158 38946 30210
rect 8766 30046 8818 30098
rect 9438 30046 9490 30098
rect 10222 30046 10274 30098
rect 15710 30046 15762 30098
rect 16606 30046 16658 30098
rect 23774 30046 23826 30098
rect 30718 30046 30770 30098
rect 35310 30046 35362 30098
rect 35534 30046 35586 30098
rect 35758 30046 35810 30098
rect 39678 30046 39730 30098
rect 14478 29934 14530 29986
rect 17614 29934 17666 29986
rect 17950 29934 18002 29986
rect 19182 29934 19234 29986
rect 20078 29934 20130 29986
rect 35086 29934 35138 29986
rect 36318 29934 36370 29986
rect 38558 29934 38610 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 16046 29598 16098 29650
rect 16718 29598 16770 29650
rect 18510 29598 18562 29650
rect 19406 29598 19458 29650
rect 30942 29598 30994 29650
rect 33518 29598 33570 29650
rect 35198 29598 35250 29650
rect 13694 29486 13746 29538
rect 15150 29486 15202 29538
rect 15934 29486 15986 29538
rect 19966 29486 20018 29538
rect 28366 29486 28418 29538
rect 34862 29486 34914 29538
rect 34974 29486 35026 29538
rect 4286 29374 4338 29426
rect 14030 29374 14082 29426
rect 14814 29374 14866 29426
rect 16270 29374 16322 29426
rect 19518 29374 19570 29426
rect 19630 29374 19682 29426
rect 19742 29374 19794 29426
rect 27694 29374 27746 29426
rect 33182 29374 33234 29426
rect 14702 29262 14754 29314
rect 17614 29262 17666 29314
rect 18062 29262 18114 29314
rect 18958 29262 19010 29314
rect 20414 29262 20466 29314
rect 24670 29262 24722 29314
rect 30494 29262 30546 29314
rect 34526 29262 34578 29314
rect 1934 29150 1986 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 14814 28814 14866 28866
rect 15486 28814 15538 28866
rect 2158 28702 2210 28754
rect 5742 28702 5794 28754
rect 7534 28702 7586 28754
rect 8990 28702 9042 28754
rect 35086 28702 35138 28754
rect 35982 28702 36034 28754
rect 39566 28702 39618 28754
rect 5070 28590 5122 28642
rect 7646 28590 7698 28642
rect 8878 28590 8930 28642
rect 9102 28590 9154 28642
rect 9326 28590 9378 28642
rect 9550 28590 9602 28642
rect 9886 28590 9938 28642
rect 14590 28590 14642 28642
rect 15150 28590 15202 28642
rect 15486 28590 15538 28642
rect 16382 28590 16434 28642
rect 16830 28590 16882 28642
rect 17838 28590 17890 28642
rect 26686 28590 26738 28642
rect 29486 28590 29538 28642
rect 4286 28478 4338 28530
rect 10446 28478 10498 28530
rect 26910 28478 26962 28530
rect 29710 28478 29762 28530
rect 34750 28478 34802 28530
rect 10110 28366 10162 28418
rect 15934 28366 15986 28418
rect 17390 28366 17442 28418
rect 34974 28366 35026 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 6302 28030 6354 28082
rect 9438 28030 9490 28082
rect 10782 28030 10834 28082
rect 14030 28030 14082 28082
rect 14142 28030 14194 28082
rect 16606 28030 16658 28082
rect 18174 28030 18226 28082
rect 22318 28030 22370 28082
rect 28590 28030 28642 28082
rect 29150 28030 29202 28082
rect 31278 28030 31330 28082
rect 32398 28030 32450 28082
rect 36318 28030 36370 28082
rect 38782 28030 38834 28082
rect 5070 27918 5122 27970
rect 8094 27918 8146 27970
rect 8990 27918 9042 27970
rect 9550 27918 9602 27970
rect 10446 27918 10498 27970
rect 14254 27918 14306 27970
rect 16382 27918 16434 27970
rect 17950 27918 18002 27970
rect 19854 27918 19906 27970
rect 20414 27918 20466 27970
rect 31502 27918 31554 27970
rect 31614 27918 31666 27970
rect 31838 27918 31890 27970
rect 32174 27918 32226 27970
rect 36654 27918 36706 27970
rect 39118 27918 39170 27970
rect 39342 27918 39394 27970
rect 39902 27918 39954 27970
rect 5742 27806 5794 27858
rect 8766 27806 8818 27858
rect 10222 27806 10274 27858
rect 11342 27806 11394 27858
rect 14814 27806 14866 27858
rect 15038 27806 15090 27858
rect 15822 27806 15874 27858
rect 17502 27806 17554 27858
rect 18398 27806 18450 27858
rect 18846 27806 18898 27858
rect 19294 27806 19346 27858
rect 20750 27806 20802 27858
rect 23102 27806 23154 27858
rect 28142 27806 28194 27858
rect 29374 27806 29426 27858
rect 33070 27806 33122 27858
rect 40238 27806 40290 27858
rect 2942 27694 2994 27746
rect 7646 27694 7698 27746
rect 7758 27694 7810 27746
rect 8206 27694 8258 27746
rect 8318 27694 8370 27746
rect 9774 27694 9826 27746
rect 9998 27694 10050 27746
rect 22766 27694 22818 27746
rect 23886 27694 23938 27746
rect 24782 27694 24834 27746
rect 25230 27694 25282 27746
rect 27358 27694 27410 27746
rect 29934 27694 29986 27746
rect 32510 27694 32562 27746
rect 33854 27694 33906 27746
rect 35982 27694 36034 27746
rect 37102 27694 37154 27746
rect 40014 27694 40066 27746
rect 8542 27582 8594 27634
rect 22318 27582 22370 27634
rect 22766 27582 22818 27634
rect 23102 27582 23154 27634
rect 23438 27582 23490 27634
rect 39454 27582 39506 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 6862 27246 6914 27298
rect 21310 27246 21362 27298
rect 22318 27246 22370 27298
rect 23998 27246 24050 27298
rect 25902 27246 25954 27298
rect 26910 27246 26962 27298
rect 2158 27134 2210 27186
rect 4286 27134 4338 27186
rect 5854 27134 5906 27186
rect 9886 27134 9938 27186
rect 11566 27134 11618 27186
rect 19966 27134 20018 27186
rect 21870 27134 21922 27186
rect 26350 27134 26402 27186
rect 27358 27134 27410 27186
rect 31950 27134 32002 27186
rect 39790 27134 39842 27186
rect 41918 27134 41970 27186
rect 5070 27022 5122 27074
rect 10446 27022 10498 27074
rect 11118 27022 11170 27074
rect 14254 27022 14306 27074
rect 14478 27022 14530 27074
rect 15822 27022 15874 27074
rect 16382 27022 16434 27074
rect 17502 27022 17554 27074
rect 18174 27022 18226 27074
rect 18398 27022 18450 27074
rect 19406 27022 19458 27074
rect 20414 27022 20466 27074
rect 21982 27022 22034 27074
rect 22318 27022 22370 27074
rect 22878 27022 22930 27074
rect 23326 27022 23378 27074
rect 23438 27022 23490 27074
rect 24110 27022 24162 27074
rect 25006 27022 25058 27074
rect 25230 27022 25282 27074
rect 25678 27022 25730 27074
rect 26238 27022 26290 27074
rect 26462 27022 26514 27074
rect 35310 27022 35362 27074
rect 35534 27022 35586 27074
rect 36318 27022 36370 27074
rect 39006 27022 39058 27074
rect 6750 26910 6802 26962
rect 10782 26910 10834 26962
rect 15934 26910 15986 26962
rect 16606 26910 16658 26962
rect 17054 26910 17106 26962
rect 19182 26910 19234 26962
rect 21422 26910 21474 26962
rect 21758 26910 21810 26962
rect 23102 26910 23154 26962
rect 25342 26910 25394 26962
rect 26798 26910 26850 26962
rect 35870 26910 35922 26962
rect 14366 26798 14418 26850
rect 16942 26798 16994 26850
rect 23662 26798 23714 26850
rect 24222 26798 24274 26850
rect 35758 26798 35810 26850
rect 38670 26798 38722 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17614 26462 17666 26514
rect 19406 26462 19458 26514
rect 19854 26462 19906 26514
rect 22542 26462 22594 26514
rect 23326 26462 23378 26514
rect 36206 26462 36258 26514
rect 7982 26350 8034 26402
rect 8878 26350 8930 26402
rect 9774 26350 9826 26402
rect 16270 26350 16322 26402
rect 19630 26350 19682 26402
rect 21534 26350 21586 26402
rect 36766 26350 36818 26402
rect 4062 26238 4114 26290
rect 8430 26238 8482 26290
rect 8654 26238 8706 26290
rect 9998 26238 10050 26290
rect 15262 26238 15314 26290
rect 15822 26238 15874 26290
rect 19966 26238 20018 26290
rect 20750 26238 20802 26290
rect 21198 26238 21250 26290
rect 21982 26238 22034 26290
rect 22878 26238 22930 26290
rect 23102 26238 23154 26290
rect 23662 26238 23714 26290
rect 24334 26238 24386 26290
rect 36542 26238 36594 26290
rect 37214 26238 37266 26290
rect 1934 26126 1986 26178
rect 8094 26126 8146 26178
rect 8206 26126 8258 26178
rect 16718 26126 16770 26178
rect 24110 26126 24162 26178
rect 25342 26126 25394 26178
rect 33182 26126 33234 26178
rect 33742 26126 33794 26178
rect 36878 26126 36930 26178
rect 37998 26126 38050 26178
rect 40238 26126 40290 26178
rect 23438 26014 23490 26066
rect 23998 26014 24050 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 6862 25678 6914 25730
rect 33518 25678 33570 25730
rect 34526 25678 34578 25730
rect 1934 25566 1986 25618
rect 14926 25566 14978 25618
rect 15710 25566 15762 25618
rect 16494 25566 16546 25618
rect 23214 25566 23266 25618
rect 29486 25566 29538 25618
rect 32846 25566 32898 25618
rect 35758 25566 35810 25618
rect 4286 25454 4338 25506
rect 14030 25454 14082 25506
rect 14702 25454 14754 25506
rect 17614 25454 17666 25506
rect 18958 25454 19010 25506
rect 19518 25454 19570 25506
rect 20414 25454 20466 25506
rect 26798 25454 26850 25506
rect 32398 25454 32450 25506
rect 33406 25454 33458 25506
rect 33630 25454 33682 25506
rect 33966 25454 34018 25506
rect 34638 25454 34690 25506
rect 35086 25454 35138 25506
rect 35310 25454 35362 25506
rect 38894 25454 38946 25506
rect 39342 25454 39394 25506
rect 39566 25454 39618 25506
rect 40126 25454 40178 25506
rect 6750 25342 6802 25394
rect 14254 25342 14306 25394
rect 14814 25342 14866 25394
rect 15038 25342 15090 25394
rect 15934 25342 15986 25394
rect 17726 25342 17778 25394
rect 19742 25342 19794 25394
rect 20302 25342 20354 25394
rect 31614 25342 31666 25394
rect 34190 25342 34242 25394
rect 34414 25342 34466 25394
rect 34862 25342 34914 25394
rect 47854 25342 47906 25394
rect 48190 25342 48242 25394
rect 15150 25230 15202 25282
rect 15710 25230 15762 25282
rect 17166 25230 17218 25282
rect 17838 25230 17890 25282
rect 18398 25230 18450 25282
rect 27246 25230 27298 25282
rect 33182 25230 33234 25282
rect 39118 25230 39170 25282
rect 47630 25230 47682 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 14814 24894 14866 24946
rect 16494 24894 16546 24946
rect 16606 24894 16658 24946
rect 17614 24894 17666 24946
rect 18510 24894 18562 24946
rect 22318 24894 22370 24946
rect 33294 24894 33346 24946
rect 34638 24894 34690 24946
rect 34974 24894 35026 24946
rect 4958 24782 5010 24834
rect 11678 24782 11730 24834
rect 13358 24782 13410 24834
rect 19854 24782 19906 24834
rect 23998 24782 24050 24834
rect 34862 24782 34914 24834
rect 36318 24782 36370 24834
rect 39118 24782 39170 24834
rect 39342 24782 39394 24834
rect 39678 24782 39730 24834
rect 5742 24670 5794 24722
rect 11790 24670 11842 24722
rect 12462 24670 12514 24722
rect 12798 24670 12850 24722
rect 16046 24670 16098 24722
rect 16382 24670 16434 24722
rect 16718 24670 16770 24722
rect 17950 24670 18002 24722
rect 18286 24670 18338 24722
rect 18398 24670 18450 24722
rect 18622 24670 18674 24722
rect 23774 24670 23826 24722
rect 30494 24670 30546 24722
rect 31054 24670 31106 24722
rect 33630 24670 33682 24722
rect 34302 24670 34354 24722
rect 36654 24670 36706 24722
rect 39454 24670 39506 24722
rect 2830 24558 2882 24610
rect 6302 24558 6354 24610
rect 11902 24558 11954 24610
rect 14590 24558 14642 24610
rect 19182 24558 19234 24610
rect 20302 24558 20354 24610
rect 27582 24558 27634 24610
rect 29710 24558 29762 24610
rect 34078 24558 34130 24610
rect 36654 24446 36706 24498
rect 39790 24446 39842 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 13022 24110 13074 24162
rect 23774 24110 23826 24162
rect 1934 23998 1986 24050
rect 7646 23998 7698 24050
rect 28590 23998 28642 24050
rect 29822 23998 29874 24050
rect 34078 23998 34130 24050
rect 36430 23998 36482 24050
rect 37774 23998 37826 24050
rect 39902 23998 39954 24050
rect 41246 23998 41298 24050
rect 43374 23998 43426 24050
rect 4286 23886 4338 23938
rect 7198 23886 7250 23938
rect 7422 23886 7474 23938
rect 7870 23886 7922 23938
rect 8206 23886 8258 23938
rect 11566 23886 11618 23938
rect 12238 23886 12290 23938
rect 12798 23886 12850 23938
rect 13918 23886 13970 23938
rect 17726 23886 17778 23938
rect 25118 23886 25170 23938
rect 29150 23886 29202 23938
rect 29486 23886 29538 23938
rect 29598 23886 29650 23938
rect 30494 23886 30546 23938
rect 30718 23886 30770 23938
rect 30830 23886 30882 23938
rect 31502 23886 31554 23938
rect 37102 23886 37154 23938
rect 40462 23886 40514 23938
rect 12686 23774 12738 23826
rect 14030 23774 14082 23826
rect 16494 23774 16546 23826
rect 23326 23774 23378 23826
rect 23662 23774 23714 23826
rect 23774 23774 23826 23826
rect 24222 23774 24274 23826
rect 24558 23774 24610 23826
rect 24894 23774 24946 23826
rect 29934 23774 29986 23826
rect 30270 23774 30322 23826
rect 7646 23662 7698 23714
rect 8542 23662 8594 23714
rect 15486 23662 15538 23714
rect 31054 23662 31106 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 24670 23326 24722 23378
rect 27582 23326 27634 23378
rect 40126 23326 40178 23378
rect 5742 23214 5794 23266
rect 7086 23214 7138 23266
rect 12686 23214 12738 23266
rect 15262 23214 15314 23266
rect 17390 23214 17442 23266
rect 20414 23214 20466 23266
rect 25566 23214 25618 23266
rect 27694 23214 27746 23266
rect 30270 23214 30322 23266
rect 4286 23102 4338 23154
rect 5854 23102 5906 23154
rect 7310 23102 7362 23154
rect 7534 23102 7586 23154
rect 7758 23102 7810 23154
rect 7982 23102 8034 23154
rect 8878 23102 8930 23154
rect 11678 23102 11730 23154
rect 12574 23102 12626 23154
rect 14702 23102 14754 23154
rect 17502 23102 17554 23154
rect 18174 23102 18226 23154
rect 18622 23102 18674 23154
rect 20302 23102 20354 23154
rect 21198 23102 21250 23154
rect 25230 23102 25282 23154
rect 27134 23102 27186 23154
rect 28254 23102 28306 23154
rect 5182 22990 5234 23042
rect 7198 22990 7250 23042
rect 8318 22990 8370 23042
rect 8654 22990 8706 23042
rect 9774 22990 9826 23042
rect 12238 22990 12290 23042
rect 13806 22990 13858 23042
rect 20750 22990 20802 23042
rect 25790 22990 25842 23042
rect 28702 22990 28754 23042
rect 29710 22990 29762 23042
rect 30382 22990 30434 23042
rect 1934 22878 1986 22930
rect 18510 22878 18562 22930
rect 27470 22878 27522 22930
rect 30046 22878 30098 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 5966 22542 6018 22594
rect 2046 22430 2098 22482
rect 4174 22430 4226 22482
rect 9886 22430 9938 22482
rect 11118 22430 11170 22482
rect 12014 22430 12066 22482
rect 14366 22430 14418 22482
rect 16382 22430 16434 22482
rect 18286 22430 18338 22482
rect 18622 22430 18674 22482
rect 21758 22430 21810 22482
rect 23774 22430 23826 22482
rect 4958 22318 5010 22370
rect 8990 22318 9042 22370
rect 10670 22318 10722 22370
rect 12574 22318 12626 22370
rect 14030 22318 14082 22370
rect 16046 22318 16098 22370
rect 29598 22318 29650 22370
rect 5854 22206 5906 22258
rect 8766 22206 8818 22258
rect 13582 22206 13634 22258
rect 14254 22206 14306 22258
rect 15150 22206 15202 22258
rect 18398 22206 18450 22258
rect 23438 22206 23490 22258
rect 24670 22206 24722 22258
rect 25230 22206 25282 22258
rect 8318 22094 8370 22146
rect 9102 22094 9154 22146
rect 9214 22094 9266 22146
rect 9326 22094 9378 22146
rect 13806 22094 13858 22146
rect 16606 22094 16658 22146
rect 20862 22094 20914 22146
rect 21310 22094 21362 22146
rect 23102 22094 23154 22146
rect 24334 22094 24386 22146
rect 24782 22094 24834 22146
rect 25006 22094 25058 22146
rect 25342 22094 25394 22146
rect 25566 22094 25618 22146
rect 25902 22094 25954 22146
rect 29822 22094 29874 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 11454 21758 11506 21810
rect 16606 21758 16658 21810
rect 19630 21758 19682 21810
rect 22206 21758 22258 21810
rect 23886 21758 23938 21810
rect 24670 21758 24722 21810
rect 34414 21758 34466 21810
rect 35198 21758 35250 21810
rect 37886 21758 37938 21810
rect 8990 21646 9042 21698
rect 10110 21646 10162 21698
rect 12574 21646 12626 21698
rect 15710 21646 15762 21698
rect 19854 21646 19906 21698
rect 20750 21646 20802 21698
rect 21534 21646 21586 21698
rect 22878 21646 22930 21698
rect 34750 21646 34802 21698
rect 4398 21534 4450 21586
rect 5182 21534 5234 21586
rect 8430 21534 8482 21586
rect 9550 21534 9602 21586
rect 9662 21534 9714 21586
rect 11566 21534 11618 21586
rect 12126 21534 12178 21586
rect 16606 21534 16658 21586
rect 19406 21534 19458 21586
rect 19966 21534 20018 21586
rect 21086 21534 21138 21586
rect 21310 21534 21362 21586
rect 21646 21534 21698 21586
rect 22542 21534 22594 21586
rect 23214 21534 23266 21586
rect 23662 21534 23714 21586
rect 2270 21422 2322 21474
rect 5630 21422 5682 21474
rect 7646 21422 7698 21474
rect 8094 21422 8146 21474
rect 14926 21422 14978 21474
rect 20526 21422 20578 21474
rect 25342 21422 25394 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 12910 20974 12962 21026
rect 22878 20974 22930 21026
rect 1934 20862 1986 20914
rect 9998 20862 10050 20914
rect 10894 20862 10946 20914
rect 12014 20862 12066 20914
rect 12350 20862 12402 20914
rect 18062 20862 18114 20914
rect 21534 20862 21586 20914
rect 24558 20862 24610 20914
rect 25566 20862 25618 20914
rect 30942 20862 30994 20914
rect 34974 20862 35026 20914
rect 41134 20862 41186 20914
rect 4286 20750 4338 20802
rect 10334 20750 10386 20802
rect 12574 20750 12626 20802
rect 14366 20750 14418 20802
rect 15374 20750 15426 20802
rect 17950 20750 18002 20802
rect 22318 20750 22370 20802
rect 22542 20750 22594 20802
rect 23774 20750 23826 20802
rect 25342 20750 25394 20802
rect 29374 20750 29426 20802
rect 29934 20750 29986 20802
rect 33854 20750 33906 20802
rect 34190 20750 34242 20802
rect 35534 20750 35586 20802
rect 37550 20750 37602 20802
rect 38222 20750 38274 20802
rect 15598 20638 15650 20690
rect 16270 20638 16322 20690
rect 20414 20638 20466 20690
rect 9102 20526 9154 20578
rect 9438 20526 9490 20578
rect 11454 20526 11506 20578
rect 13806 20526 13858 20578
rect 21982 20526 22034 20578
rect 23214 20526 23266 20578
rect 25006 20526 25058 20578
rect 25902 20526 25954 20578
rect 28590 20526 28642 20578
rect 29598 20526 29650 20578
rect 29710 20582 29762 20634
rect 30158 20638 30210 20690
rect 30382 20638 30434 20690
rect 30606 20638 30658 20690
rect 33070 20638 33122 20690
rect 36990 20638 37042 20690
rect 37214 20638 37266 20690
rect 37438 20638 37490 20690
rect 39006 20638 39058 20690
rect 34526 20526 34578 20578
rect 35758 20526 35810 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 12238 20190 12290 20242
rect 24222 20190 24274 20242
rect 30494 20190 30546 20242
rect 2046 20078 2098 20130
rect 8990 20078 9042 20130
rect 10110 20078 10162 20130
rect 11678 20078 11730 20130
rect 12910 20078 12962 20130
rect 14702 20078 14754 20130
rect 15374 20078 15426 20130
rect 24670 20078 24722 20130
rect 26350 20078 26402 20130
rect 26462 20078 26514 20130
rect 27022 20078 27074 20130
rect 30718 20078 30770 20130
rect 31838 20078 31890 20130
rect 34526 20078 34578 20130
rect 34974 20078 35026 20130
rect 35534 20078 35586 20130
rect 35758 20078 35810 20130
rect 47854 20078 47906 20130
rect 1710 19966 1762 20018
rect 8766 19966 8818 20018
rect 12798 19966 12850 20018
rect 16606 19966 16658 20018
rect 20750 19966 20802 20018
rect 21310 19966 21362 20018
rect 25454 19966 25506 20018
rect 25678 19966 25730 20018
rect 26686 19966 26738 20018
rect 30830 19966 30882 20018
rect 32062 19966 32114 20018
rect 34862 19966 34914 20018
rect 35198 19966 35250 20018
rect 35422 19966 35474 20018
rect 36318 19966 36370 20018
rect 36542 19966 36594 20018
rect 36766 19966 36818 20018
rect 37326 19966 37378 20018
rect 48190 19966 48242 20018
rect 2494 19854 2546 19906
rect 7982 19854 8034 19906
rect 8318 19854 8370 19906
rect 9774 19854 9826 19906
rect 10670 19854 10722 19906
rect 11006 19854 11058 19906
rect 11342 19854 11394 19906
rect 11902 19854 11954 19906
rect 20414 19854 20466 19906
rect 22878 19854 22930 19906
rect 23326 19854 23378 19906
rect 30270 19854 30322 19906
rect 36430 19854 36482 19906
rect 37998 19854 38050 19906
rect 40126 19854 40178 19906
rect 47630 19854 47682 19906
rect 22878 19742 22930 19794
rect 23214 19742 23266 19794
rect 26014 19742 26066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 11566 19406 11618 19458
rect 12462 19406 12514 19458
rect 14030 19406 14082 19458
rect 14366 19406 14418 19458
rect 15934 19406 15986 19458
rect 36318 19406 36370 19458
rect 37102 19406 37154 19458
rect 10670 19294 10722 19346
rect 12350 19294 12402 19346
rect 13806 19294 13858 19346
rect 16158 19294 16210 19346
rect 16718 19294 16770 19346
rect 19966 19294 20018 19346
rect 27918 19294 27970 19346
rect 35198 19294 35250 19346
rect 37662 19294 37714 19346
rect 38110 19294 38162 19346
rect 9774 19182 9826 19234
rect 11006 19182 11058 19234
rect 12014 19182 12066 19234
rect 12126 19182 12178 19234
rect 15262 19182 15314 19234
rect 26798 19182 26850 19234
rect 30606 19182 30658 19234
rect 31950 19182 32002 19234
rect 36430 19182 36482 19234
rect 36990 19182 37042 19234
rect 15150 19070 15202 19122
rect 19406 19070 19458 19122
rect 19518 19070 19570 19122
rect 27246 19070 27298 19122
rect 27470 19070 27522 19122
rect 31278 19070 31330 19122
rect 31726 19070 31778 19122
rect 37102 19070 37154 19122
rect 8878 18958 8930 19010
rect 9214 18958 9266 19010
rect 10110 18958 10162 19010
rect 14926 18958 14978 19010
rect 15598 18958 15650 19010
rect 18174 18958 18226 19010
rect 19182 18958 19234 19010
rect 27134 18958 27186 19010
rect 29262 18958 29314 19010
rect 30718 18958 30770 19010
rect 30942 18958 30994 19010
rect 32734 18958 32786 19010
rect 35870 18958 35922 19010
rect 36318 18958 36370 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 11118 18622 11170 18674
rect 15150 18622 15202 18674
rect 16270 18622 16322 18674
rect 25678 18622 25730 18674
rect 2046 18510 2098 18562
rect 9774 18510 9826 18562
rect 11566 18510 11618 18562
rect 13022 18510 13074 18562
rect 15598 18510 15650 18562
rect 18062 18510 18114 18562
rect 18174 18510 18226 18562
rect 27918 18510 27970 18562
rect 29374 18510 29426 18562
rect 37662 18510 37714 18562
rect 1710 18398 1762 18450
rect 6526 18398 6578 18450
rect 7198 18398 7250 18450
rect 11902 18398 11954 18450
rect 13918 18398 13970 18450
rect 18510 18398 18562 18450
rect 24110 18398 24162 18450
rect 28702 18398 28754 18450
rect 29038 18398 29090 18450
rect 30494 18398 30546 18450
rect 32174 18398 32226 18450
rect 33294 18398 33346 18450
rect 2494 18286 2546 18338
rect 6638 18286 6690 18338
rect 7646 18286 7698 18338
rect 8094 18286 8146 18338
rect 10670 18286 10722 18338
rect 17614 18286 17666 18338
rect 19294 18286 19346 18338
rect 21422 18286 21474 18338
rect 23774 18286 23826 18338
rect 24558 18286 24610 18338
rect 29822 18286 29874 18338
rect 31390 18286 31442 18338
rect 31838 18286 31890 18338
rect 32510 18286 32562 18338
rect 6078 18174 6130 18226
rect 7198 18174 7250 18226
rect 7646 18174 7698 18226
rect 8206 18174 8258 18226
rect 18062 18174 18114 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 30158 17838 30210 17890
rect 5070 17726 5122 17778
rect 8094 17726 8146 17778
rect 9774 17726 9826 17778
rect 19406 17726 19458 17778
rect 20750 17726 20802 17778
rect 25342 17726 25394 17778
rect 25678 17726 25730 17778
rect 27022 17726 27074 17778
rect 32846 17726 32898 17778
rect 2270 17614 2322 17666
rect 7198 17614 7250 17666
rect 7870 17614 7922 17666
rect 18398 17614 18450 17666
rect 19182 17614 19234 17666
rect 19518 17614 19570 17666
rect 19742 17614 19794 17666
rect 26126 17614 26178 17666
rect 27246 17614 27298 17666
rect 29486 17614 29538 17666
rect 29934 17614 29986 17666
rect 31278 17614 31330 17666
rect 31614 17614 31666 17666
rect 35982 17614 36034 17666
rect 2942 17502 2994 17554
rect 6078 17502 6130 17554
rect 6190 17502 6242 17554
rect 6414 17502 6466 17554
rect 6638 17502 6690 17554
rect 6750 17502 6802 17554
rect 6974 17502 7026 17554
rect 8206 17502 8258 17554
rect 8430 17502 8482 17554
rect 8654 17502 8706 17554
rect 8766 17502 8818 17554
rect 9214 17502 9266 17554
rect 9326 17502 9378 17554
rect 15038 17502 15090 17554
rect 20302 17502 20354 17554
rect 27470 17502 27522 17554
rect 27582 17502 27634 17554
rect 30606 17502 30658 17554
rect 30718 17502 30770 17554
rect 31950 17502 32002 17554
rect 5742 17390 5794 17442
rect 8990 17390 9042 17442
rect 28254 17390 28306 17442
rect 28590 17390 28642 17442
rect 30942 17390 30994 17442
rect 31614 17390 31666 17442
rect 36094 17390 36146 17442
rect 36318 17390 36370 17442
rect 37102 17390 37154 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 7758 17054 7810 17106
rect 8542 17054 8594 17106
rect 9102 17054 9154 17106
rect 11006 17054 11058 17106
rect 18622 17054 18674 17106
rect 19406 17054 19458 17106
rect 19854 17054 19906 17106
rect 21310 17054 21362 17106
rect 29150 17054 29202 17106
rect 30382 17054 30434 17106
rect 30942 17054 30994 17106
rect 31166 17054 31218 17106
rect 31502 17054 31554 17106
rect 33742 17054 33794 17106
rect 37662 17054 37714 17106
rect 4062 16942 4114 16994
rect 6750 16942 6802 16994
rect 6862 16942 6914 16994
rect 7086 16942 7138 16994
rect 7534 16942 7586 16994
rect 10670 16942 10722 16994
rect 18958 16942 19010 16994
rect 19742 16942 19794 16994
rect 20078 16942 20130 16994
rect 20302 16942 20354 16994
rect 20750 16942 20802 16994
rect 20862 16942 20914 16994
rect 22542 16942 22594 16994
rect 30830 16942 30882 16994
rect 33182 16942 33234 16994
rect 35534 16942 35586 16994
rect 36206 16942 36258 16994
rect 1822 16830 1874 16882
rect 2270 16830 2322 16882
rect 3390 16830 3442 16882
rect 7198 16830 7250 16882
rect 7870 16830 7922 16882
rect 20638 16830 20690 16882
rect 21086 16830 21138 16882
rect 21422 16830 21474 16882
rect 21870 16830 21922 16882
rect 25454 16830 25506 16882
rect 33070 16830 33122 16882
rect 33406 16830 33458 16882
rect 35422 16830 35474 16882
rect 35982 16830 36034 16882
rect 36430 16830 36482 16882
rect 36654 16830 36706 16882
rect 37214 16830 37266 16882
rect 6190 16718 6242 16770
rect 24670 16718 24722 16770
rect 35758 16718 35810 16770
rect 36318 16718 36370 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 35982 16270 36034 16322
rect 1822 16158 1874 16210
rect 5742 16158 5794 16210
rect 14366 16158 14418 16210
rect 16158 16158 16210 16210
rect 17054 16158 17106 16210
rect 17950 16158 18002 16210
rect 20078 16158 20130 16210
rect 21646 16158 21698 16210
rect 32734 16158 32786 16210
rect 34862 16158 34914 16210
rect 35534 16158 35586 16210
rect 37774 16158 37826 16210
rect 40014 16158 40066 16210
rect 6078 16046 6130 16098
rect 6974 16046 7026 16098
rect 7198 16046 7250 16098
rect 7870 16046 7922 16098
rect 8206 16046 8258 16098
rect 9998 16046 10050 16098
rect 12910 16046 12962 16098
rect 13806 16046 13858 16098
rect 17390 16046 17442 16098
rect 31726 16046 31778 16098
rect 32062 16046 32114 16098
rect 36094 16046 36146 16098
rect 36990 16046 37042 16098
rect 6190 15934 6242 15986
rect 6414 15934 6466 15986
rect 6638 15934 6690 15986
rect 8094 15934 8146 15986
rect 8654 15934 8706 15986
rect 9774 15934 9826 15986
rect 14702 15934 14754 15986
rect 14814 15934 14866 15986
rect 15262 15934 15314 15986
rect 15374 15934 15426 15986
rect 31390 15934 31442 15986
rect 31502 15934 31554 15986
rect 5182 15822 5234 15874
rect 6750 15822 6802 15874
rect 7646 15822 7698 15874
rect 13470 15822 13522 15874
rect 15038 15822 15090 15874
rect 15598 15822 15650 15874
rect 16494 15822 16546 15874
rect 20638 15822 20690 15874
rect 20862 15822 20914 15874
rect 31166 15822 31218 15874
rect 35982 15822 36034 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 6862 15486 6914 15538
rect 7422 15486 7474 15538
rect 7758 15486 7810 15538
rect 9550 15486 9602 15538
rect 12462 15486 12514 15538
rect 12798 15486 12850 15538
rect 13246 15486 13298 15538
rect 17502 15486 17554 15538
rect 19854 15486 19906 15538
rect 20302 15486 20354 15538
rect 20638 15486 20690 15538
rect 26014 15486 26066 15538
rect 29934 15486 29986 15538
rect 30270 15486 30322 15538
rect 31726 15486 31778 15538
rect 31950 15486 32002 15538
rect 39902 15486 39954 15538
rect 3166 15374 3218 15426
rect 6190 15374 6242 15426
rect 10334 15374 10386 15426
rect 10446 15374 10498 15426
rect 13134 15374 13186 15426
rect 19742 15374 19794 15426
rect 21646 15374 21698 15426
rect 21982 15374 22034 15426
rect 22094 15374 22146 15426
rect 37102 15374 37154 15426
rect 2494 15262 2546 15314
rect 6302 15262 6354 15314
rect 9886 15262 9938 15314
rect 10110 15262 10162 15314
rect 14030 15262 14082 15314
rect 20974 15262 21026 15314
rect 21422 15262 21474 15314
rect 22318 15262 22370 15314
rect 22654 15262 22706 15314
rect 26798 15262 26850 15314
rect 28590 15262 28642 15314
rect 30158 15262 30210 15314
rect 30494 15262 30546 15314
rect 36318 15262 36370 15314
rect 1822 15150 1874 15202
rect 5294 15150 5346 15202
rect 5630 15150 5682 15202
rect 10894 15150 10946 15202
rect 14702 15150 14754 15202
rect 16830 15150 16882 15202
rect 19406 15150 19458 15202
rect 21198 15150 21250 15202
rect 26462 15150 26514 15202
rect 32398 15150 32450 15202
rect 39230 15150 39282 15202
rect 13246 15038 13298 15090
rect 19854 15038 19906 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19966 14702 20018 14754
rect 5854 14590 5906 14642
rect 6302 14590 6354 14642
rect 12014 14590 12066 14642
rect 14814 14590 14866 14642
rect 18286 14590 18338 14642
rect 27134 14590 27186 14642
rect 1710 14478 1762 14530
rect 2270 14478 2322 14530
rect 9326 14478 9378 14530
rect 11006 14478 11058 14530
rect 12574 14478 12626 14530
rect 14366 14478 14418 14530
rect 14590 14478 14642 14530
rect 15038 14478 15090 14530
rect 18846 14478 18898 14530
rect 19854 14478 19906 14530
rect 21198 14478 21250 14530
rect 21646 14478 21698 14530
rect 21870 14478 21922 14530
rect 26126 14478 26178 14530
rect 27582 14478 27634 14530
rect 28030 14478 28082 14530
rect 30158 14478 30210 14530
rect 12462 14366 12514 14418
rect 15262 14366 15314 14418
rect 16270 14366 16322 14418
rect 18734 14366 18786 14418
rect 8990 14254 9042 14306
rect 9438 14254 9490 14306
rect 9662 14254 9714 14306
rect 11230 14254 11282 14306
rect 12238 14254 12290 14306
rect 13918 14254 13970 14306
rect 14030 14254 14082 14306
rect 14254 14254 14306 14306
rect 15934 14254 15986 14306
rect 18510 14254 18562 14306
rect 19630 14254 19682 14306
rect 19966 14254 20018 14306
rect 20414 14310 20466 14362
rect 28366 14366 28418 14418
rect 32062 14366 32114 14418
rect 48190 14366 48242 14418
rect 20526 14254 20578 14306
rect 20750 14254 20802 14306
rect 21422 14254 21474 14306
rect 25678 14254 25730 14306
rect 26350 14254 26402 14306
rect 26686 14254 26738 14306
rect 47630 14254 47682 14306
rect 47854 14254 47906 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 11454 13918 11506 13970
rect 27246 13918 27298 13970
rect 27918 13918 27970 13970
rect 28926 13918 28978 13970
rect 29374 13918 29426 13970
rect 9550 13806 9602 13858
rect 9886 13806 9938 13858
rect 10446 13806 10498 13858
rect 10782 13806 10834 13858
rect 22542 13806 22594 13858
rect 28030 13806 28082 13858
rect 28478 13806 28530 13858
rect 29822 13806 29874 13858
rect 30046 13806 30098 13858
rect 30270 13806 30322 13858
rect 30830 13806 30882 13858
rect 1822 13694 1874 13746
rect 2270 13694 2322 13746
rect 10110 13694 10162 13746
rect 20862 13694 20914 13746
rect 21758 13694 21810 13746
rect 27694 13694 27746 13746
rect 29710 13694 29762 13746
rect 30494 13694 30546 13746
rect 31054 13694 31106 13746
rect 31390 13694 31442 13746
rect 31614 13694 31666 13746
rect 9662 13582 9714 13634
rect 21534 13582 21586 13634
rect 24670 13582 24722 13634
rect 30382 13582 30434 13634
rect 31278 13582 31330 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 1822 13022 1874 13074
rect 20302 13022 20354 13074
rect 24222 13022 24274 13074
rect 26350 13022 26402 13074
rect 28590 13022 28642 13074
rect 32734 13022 32786 13074
rect 34862 13022 34914 13074
rect 11454 12910 11506 12962
rect 11678 12910 11730 12962
rect 12686 12910 12738 12962
rect 13022 12910 13074 12962
rect 13358 12910 13410 12962
rect 13694 12910 13746 12962
rect 13918 12910 13970 12962
rect 14590 12910 14642 12962
rect 16718 12910 16770 12962
rect 21534 12910 21586 12962
rect 23550 12910 23602 12962
rect 27806 12910 27858 12962
rect 29262 12910 29314 12962
rect 30046 12910 30098 12962
rect 30718 12910 30770 12962
rect 32062 12910 32114 12962
rect 11902 12798 11954 12850
rect 14478 12798 14530 12850
rect 27246 12798 27298 12850
rect 29374 12798 29426 12850
rect 30382 12798 30434 12850
rect 11790 12686 11842 12738
rect 12462 12686 12514 12738
rect 12798 12686 12850 12738
rect 13582 12686 13634 12738
rect 14254 12686 14306 12738
rect 26798 12686 26850 12738
rect 27470 12686 27522 12738
rect 27694 12686 27746 12738
rect 29598 12686 29650 12738
rect 29710 12686 29762 12738
rect 29934 12686 29986 12738
rect 30494 12686 30546 12738
rect 31054 12686 31106 12738
rect 31502 12686 31554 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 11678 12350 11730 12402
rect 11902 12350 11954 12402
rect 12126 12350 12178 12402
rect 14814 12350 14866 12402
rect 27694 12350 27746 12402
rect 8206 12238 8258 12290
rect 12238 12238 12290 12290
rect 13358 12238 13410 12290
rect 13582 12238 13634 12290
rect 18958 12238 19010 12290
rect 20526 12238 20578 12290
rect 27470 12238 27522 12290
rect 29822 12238 29874 12290
rect 1822 12126 1874 12178
rect 8990 12126 9042 12178
rect 14030 12126 14082 12178
rect 18846 12126 18898 12178
rect 19294 12126 19346 12178
rect 20750 12126 20802 12178
rect 27694 12126 27746 12178
rect 27918 12126 27970 12178
rect 28590 12126 28642 12178
rect 29262 12126 29314 12178
rect 29598 12126 29650 12178
rect 30382 12126 30434 12178
rect 2270 12014 2322 12066
rect 6078 12014 6130 12066
rect 9662 12014 9714 12066
rect 13806 12014 13858 12066
rect 19182 12014 19234 12066
rect 29710 12014 29762 12066
rect 31614 12014 31666 12066
rect 28142 11902 28194 11954
rect 28478 11902 28530 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 21646 11566 21698 11618
rect 1822 11454 1874 11506
rect 14814 11454 14866 11506
rect 16494 11454 16546 11506
rect 18062 11454 18114 11506
rect 20190 11454 20242 11506
rect 21982 11454 22034 11506
rect 33966 11454 34018 11506
rect 15598 11342 15650 11394
rect 15822 11342 15874 11394
rect 16942 11342 16994 11394
rect 17390 11342 17442 11394
rect 20750 11342 20802 11394
rect 30942 11342 30994 11394
rect 31726 11342 31778 11394
rect 15934 11230 15986 11282
rect 21870 11230 21922 11282
rect 34526 11118 34578 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 14926 10782 14978 10834
rect 16494 10782 16546 10834
rect 19182 10782 19234 10834
rect 20078 10782 20130 10834
rect 20638 10782 20690 10834
rect 20974 10782 21026 10834
rect 26238 10782 26290 10834
rect 2270 10670 2322 10722
rect 13694 10670 13746 10722
rect 19406 10670 19458 10722
rect 21198 10670 21250 10722
rect 21870 10670 21922 10722
rect 28478 10670 28530 10722
rect 1822 10558 1874 10610
rect 14478 10558 14530 10610
rect 15374 10558 15426 10610
rect 15822 10558 15874 10610
rect 19518 10558 19570 10610
rect 21646 10558 21698 10610
rect 29150 10558 29202 10610
rect 11566 10446 11618 10498
rect 29710 10446 29762 10498
rect 15374 10334 15426 10386
rect 20862 10334 20914 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 20302 9998 20354 10050
rect 22318 9998 22370 10050
rect 1822 9886 1874 9938
rect 9438 9886 9490 9938
rect 11566 9886 11618 9938
rect 12126 9886 12178 9938
rect 15374 9886 15426 9938
rect 19966 9886 20018 9938
rect 23102 9886 23154 9938
rect 29934 9886 29986 9938
rect 32734 9886 32786 9938
rect 8766 9774 8818 9826
rect 12462 9774 12514 9826
rect 14142 9774 14194 9826
rect 14366 9774 14418 9826
rect 15710 9774 15762 9826
rect 21870 9774 21922 9826
rect 22206 9774 22258 9826
rect 22430 9774 22482 9826
rect 23550 9774 23602 9826
rect 24334 9774 24386 9826
rect 29150 9774 29202 9826
rect 13582 9662 13634 9714
rect 24446 9662 24498 9714
rect 12574 9550 12626 9602
rect 14814 9550 14866 9602
rect 19630 9550 19682 9602
rect 20078 9550 20130 9602
rect 22654 9550 22706 9602
rect 32174 9550 32226 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 2046 9214 2098 9266
rect 11454 9214 11506 9266
rect 11790 9214 11842 9266
rect 12350 9214 12402 9266
rect 15934 9214 15986 9266
rect 18622 9214 18674 9266
rect 20078 9214 20130 9266
rect 13358 9102 13410 9154
rect 19518 9102 19570 9154
rect 20190 9102 20242 9154
rect 20526 9102 20578 9154
rect 20750 9102 20802 9154
rect 22206 9102 22258 9154
rect 47854 9102 47906 9154
rect 1710 8990 1762 9042
rect 12686 8990 12738 9042
rect 19182 8990 19234 9042
rect 19294 8990 19346 9042
rect 19742 8990 19794 9042
rect 20974 8990 21026 9042
rect 21310 8990 21362 9042
rect 25902 8990 25954 9042
rect 26238 8990 26290 9042
rect 48190 8990 48242 9042
rect 2494 8878 2546 8930
rect 15486 8878 15538 8930
rect 19630 8878 19682 8930
rect 20638 8878 20690 8930
rect 21758 8878 21810 8930
rect 26686 8878 26738 8930
rect 27134 8878 27186 8930
rect 47630 8878 47682 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 20078 8318 20130 8370
rect 23662 8318 23714 8370
rect 25790 8318 25842 8370
rect 22990 8206 23042 8258
rect 26350 8206 26402 8258
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 2046 7646 2098 7698
rect 16830 7646 16882 7698
rect 21870 7646 21922 7698
rect 19518 7534 19570 7586
rect 1710 7422 1762 7474
rect 20190 7422 20242 7474
rect 20638 7422 20690 7474
rect 21086 7422 21138 7474
rect 2494 7310 2546 7362
rect 17390 7310 17442 7362
rect 21310 7198 21362 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 22654 6862 22706 6914
rect 23438 6862 23490 6914
rect 20414 6750 20466 6802
rect 22430 6750 22482 6802
rect 23662 6638 23714 6690
rect 24222 6638 24274 6690
rect 22766 6526 22818 6578
rect 23102 6414 23154 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 19742 6078 19794 6130
rect 20862 5966 20914 6018
rect 1822 5854 1874 5906
rect 2270 5854 2322 5906
rect 20190 5854 20242 5906
rect 22990 5742 23042 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 1822 5182 1874 5234
rect 24110 5182 24162 5234
rect 22542 5070 22594 5122
rect 23102 5070 23154 5122
rect 22766 4958 22818 5010
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 2046 4510 2098 4562
rect 22094 4510 22146 4562
rect 40350 4510 40402 4562
rect 47854 4510 47906 4562
rect 1710 4286 1762 4338
rect 7086 4286 7138 4338
rect 12014 4286 12066 4338
rect 13358 4286 13410 4338
rect 21646 4286 21698 4338
rect 27134 4286 27186 4338
rect 33182 4286 33234 4338
rect 41246 4286 41298 4338
rect 48190 4286 48242 4338
rect 2494 4174 2546 4226
rect 2942 4174 2994 4226
rect 46958 4174 47010 4226
rect 47630 4174 47682 4226
rect 5182 4062 5234 4114
rect 9774 4062 9826 4114
rect 14030 4062 14082 4114
rect 19294 4062 19346 4114
rect 28142 4062 28194 4114
rect 34190 4062 34242 4114
rect 42254 4062 42306 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 2718 3614 2770 3666
rect 6750 3614 6802 3666
rect 17278 3614 17330 3666
rect 22094 3614 22146 3666
rect 25342 3614 25394 3666
rect 40014 3614 40066 3666
rect 42814 3614 42866 3666
rect 43822 3614 43874 3666
rect 47854 3614 47906 3666
rect 4958 3502 5010 3554
rect 8318 3502 8370 3554
rect 12574 3502 12626 3554
rect 16046 3502 16098 3554
rect 19182 3502 19234 3554
rect 20078 3502 20130 3554
rect 21310 3502 21362 3554
rect 27246 3502 27298 3554
rect 28478 3502 28530 3554
rect 29038 3502 29090 3554
rect 32622 3502 32674 3554
rect 36206 3502 36258 3554
rect 37438 3502 37490 3554
rect 42030 3502 42082 3554
rect 45726 3502 45778 3554
rect 46622 3502 46674 3554
rect 1710 3390 1762 3442
rect 2046 3390 2098 3442
rect 10782 3390 10834 3442
rect 14814 3390 14866 3442
rect 33742 3390 33794 3442
rect 35534 3390 35586 3442
rect 35982 3390 36034 3442
rect 36990 3390 37042 3442
rect 37214 3390 37266 3442
rect 47406 3390 47458 3442
rect 30046 3278 30098 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 2688 49200 2800 50000
rect 4032 49200 4144 50000
rect 5376 49200 5488 50000
rect 6720 49200 6832 50000
rect 8064 49200 8176 50000
rect 9408 49200 9520 50000
rect 10752 49200 10864 50000
rect 12096 49200 12208 50000
rect 13440 49200 13552 50000
rect 14784 49200 14896 50000
rect 16128 49200 16240 50000
rect 17472 49200 17584 50000
rect 18816 49200 18928 50000
rect 20160 49200 20272 50000
rect 21504 49200 21616 50000
rect 22848 49200 22960 50000
rect 24192 49200 24304 50000
rect 25536 49200 25648 50000
rect 25900 49308 26292 49364
rect 2716 46900 2772 49200
rect 2716 46834 2772 46844
rect 1932 46004 1988 46014
rect 1932 45910 1988 45948
rect 3948 45106 4004 45118
rect 3948 45054 3950 45106
rect 4002 45054 4004 45106
rect 1932 44884 1988 44894
rect 1820 44882 1988 44884
rect 1820 44830 1934 44882
rect 1986 44830 1988 44882
rect 1820 44828 1988 44830
rect 1820 44436 1876 44828
rect 1932 44818 1988 44828
rect 1820 44370 1876 44380
rect 1932 44434 1988 44446
rect 1932 44382 1934 44434
rect 1986 44382 1988 44434
rect 1596 44324 1652 44334
rect 1484 43876 1540 43886
rect 1484 29876 1540 43820
rect 1484 29810 1540 29820
rect 1596 26516 1652 44268
rect 1932 43708 1988 44382
rect 1932 43652 2212 43708
rect 1932 43314 1988 43326
rect 1932 43262 1934 43314
rect 1986 43262 1988 43314
rect 1932 42868 1988 43262
rect 1932 42802 1988 42812
rect 2044 42866 2100 42878
rect 2044 42814 2046 42866
rect 2098 42814 2100 42866
rect 2044 41412 2100 42814
rect 2044 41346 2100 41356
rect 2156 42868 2212 43652
rect 2044 41186 2100 41198
rect 2044 41134 2046 41186
rect 2098 41134 2100 41186
rect 2044 40964 2100 41134
rect 2044 40898 2100 40908
rect 1932 40178 1988 40190
rect 1932 40126 1934 40178
rect 1986 40126 1988 40178
rect 1932 39732 1988 40126
rect 1932 39666 1988 39676
rect 1932 38610 1988 38622
rect 1932 38558 1934 38610
rect 1986 38558 1988 38610
rect 1932 38164 1988 38558
rect 1932 38098 1988 38108
rect 2156 38164 2212 42812
rect 3948 42644 4004 45054
rect 4060 44436 4116 49200
rect 4844 47572 4900 47582
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4284 45890 4340 45902
rect 4284 45838 4286 45890
rect 4338 45838 4340 45890
rect 4284 45556 4340 45838
rect 4732 45892 4788 45902
rect 4732 45798 4788 45836
rect 4284 45490 4340 45500
rect 4844 44994 4900 47516
rect 5404 45892 5460 49200
rect 4844 44942 4846 44994
rect 4898 44942 4900 44994
rect 4844 44930 4900 44942
rect 4956 45666 5012 45678
rect 4956 45614 4958 45666
rect 5010 45614 5012 45666
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4060 44380 4788 44436
rect 3948 42578 4004 42588
rect 4060 44210 4116 44222
rect 4060 44158 4062 44210
rect 4114 44158 4116 44210
rect 3836 41970 3892 41982
rect 3836 41918 3838 41970
rect 3890 41918 3892 41970
rect 2716 41074 2772 41086
rect 2716 41022 2718 41074
rect 2770 41022 2772 41074
rect 2716 39508 2772 41022
rect 3836 40964 3892 41918
rect 3836 40898 3892 40908
rect 2716 39452 3444 39508
rect 2156 38098 2212 38108
rect 2828 38164 2884 38174
rect 2828 38070 2884 38108
rect 3388 38162 3444 39452
rect 3836 38724 3892 38734
rect 3836 38276 3892 38668
rect 3388 38110 3390 38162
rect 3442 38110 3444 38162
rect 3388 38098 3444 38110
rect 3500 38220 3892 38276
rect 3276 38052 3332 38062
rect 3276 37958 3332 37996
rect 3500 37940 3556 38220
rect 3388 37884 3556 37940
rect 3612 38050 3668 38062
rect 3612 37998 3614 38050
rect 3666 37998 3668 38050
rect 2940 37826 2996 37838
rect 2940 37774 2942 37826
rect 2994 37774 2996 37826
rect 2380 37268 2436 37278
rect 2380 37174 2436 37212
rect 2940 36708 2996 37774
rect 2940 36642 2996 36652
rect 3052 37154 3108 37166
rect 3052 37102 3054 37154
rect 3106 37102 3108 37154
rect 1932 36596 1988 36606
rect 1932 36502 1988 36540
rect 3052 35924 3108 37102
rect 3052 35858 3108 35868
rect 1932 35474 1988 35486
rect 1932 35422 1934 35474
rect 1986 35422 1988 35474
rect 1932 35028 1988 35422
rect 1932 34962 1988 34972
rect 2044 35476 2100 35486
rect 2044 34354 2100 35420
rect 3388 35364 3444 37884
rect 3612 37604 3668 37998
rect 3612 37538 3668 37548
rect 3724 38050 3780 38062
rect 3724 37998 3726 38050
rect 3778 37998 3780 38050
rect 3276 35308 3444 35364
rect 3500 35924 3556 35934
rect 3164 35028 3220 35038
rect 2828 34916 2884 34926
rect 2828 34822 2884 34860
rect 2940 34804 2996 34814
rect 2940 34710 2996 34748
rect 2380 34692 2436 34702
rect 2716 34692 2772 34702
rect 2380 34690 2772 34692
rect 2380 34638 2382 34690
rect 2434 34638 2718 34690
rect 2770 34638 2772 34690
rect 2380 34636 2772 34638
rect 2380 34626 2436 34636
rect 2044 34302 2046 34354
rect 2098 34302 2100 34354
rect 2044 34290 2100 34302
rect 2716 34244 2772 34636
rect 2716 34178 2772 34188
rect 3052 34244 3108 34254
rect 1708 34130 1764 34142
rect 1708 34078 1710 34130
rect 1762 34078 1764 34130
rect 1708 33460 1764 34078
rect 1708 33394 1764 33404
rect 2492 34018 2548 34030
rect 2492 33966 2494 34018
rect 2546 33966 2548 34018
rect 2492 33460 2548 33966
rect 2492 33394 2548 33404
rect 1932 32340 1988 32350
rect 1820 32338 1988 32340
rect 1820 32286 1934 32338
rect 1986 32286 1988 32338
rect 1820 32284 1988 32286
rect 1820 31892 1876 32284
rect 1932 32274 1988 32284
rect 1820 31826 1876 31836
rect 1932 31890 1988 31902
rect 1932 31838 1934 31890
rect 1986 31838 1988 31890
rect 1932 31780 1988 31838
rect 1932 31714 1988 31724
rect 1932 30324 1988 30334
rect 1932 30230 1988 30268
rect 1932 29202 1988 29214
rect 1932 29150 1934 29202
rect 1986 29150 1988 29202
rect 1932 28756 1988 29150
rect 1932 28690 1988 28700
rect 2156 28756 2212 28766
rect 2156 28662 2212 28700
rect 2940 27746 2996 27758
rect 2940 27694 2942 27746
rect 2994 27694 2996 27746
rect 2940 27636 2996 27694
rect 2940 27570 2996 27580
rect 1596 26450 1652 26460
rect 1932 27188 1988 27198
rect 1932 26178 1988 27132
rect 2156 27186 2212 27198
rect 2156 27134 2158 27186
rect 2210 27134 2212 27186
rect 2156 26964 2212 27134
rect 2156 26898 2212 26908
rect 1932 26126 1934 26178
rect 1986 26126 1988 26178
rect 1932 26114 1988 26126
rect 1932 25620 1988 25630
rect 1932 25526 1988 25564
rect 2828 24612 2884 24622
rect 2828 24518 2884 24556
rect 1932 24052 1988 24062
rect 1932 23958 1988 23996
rect 2044 23156 2100 23166
rect 1932 22930 1988 22942
rect 1932 22878 1934 22930
rect 1986 22878 1988 22930
rect 1932 22484 1988 22878
rect 1932 22418 1988 22428
rect 2044 22482 2100 23100
rect 2044 22430 2046 22482
rect 2098 22430 2100 22482
rect 2044 22418 2100 22430
rect 2268 21474 2324 21486
rect 2268 21422 2270 21474
rect 2322 21422 2324 21474
rect 1932 20916 1988 20926
rect 1932 20822 1988 20860
rect 2268 20804 2324 21422
rect 2268 20738 2324 20748
rect 2044 20130 2100 20142
rect 2044 20078 2046 20130
rect 2098 20078 2100 20130
rect 1708 20018 1764 20030
rect 1708 19966 1710 20018
rect 1762 19966 1764 20018
rect 1708 19908 1764 19966
rect 1708 19348 1764 19852
rect 2044 19796 2100 20078
rect 2492 19908 2548 19918
rect 2492 19814 2548 19852
rect 2044 19730 2100 19740
rect 1708 19282 1764 19292
rect 1932 19124 1988 19134
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18340 1764 18398
rect 1708 17780 1764 18284
rect 1708 17714 1764 17724
rect 1820 16882 1876 16894
rect 1820 16830 1822 16882
rect 1874 16830 1876 16882
rect 1820 16212 1876 16830
rect 1820 16118 1876 16156
rect 1820 15202 1876 15214
rect 1820 15150 1822 15202
rect 1874 15150 1876 15202
rect 1708 14644 1764 14654
rect 1820 14644 1876 15150
rect 1764 14588 1876 14644
rect 1708 14530 1764 14588
rect 1708 14478 1710 14530
rect 1762 14478 1764 14530
rect 1708 14466 1764 14478
rect 1820 13746 1876 13758
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 13076 1876 13694
rect 1820 12982 1876 13020
rect 1820 12178 1876 12190
rect 1820 12126 1822 12178
rect 1874 12126 1876 12178
rect 1820 11508 1876 12126
rect 1820 11414 1876 11452
rect 1820 10610 1876 10622
rect 1820 10558 1822 10610
rect 1874 10558 1876 10610
rect 1820 9940 1876 10558
rect 1820 9846 1876 9884
rect 1708 9042 1764 9054
rect 1708 8990 1710 9042
rect 1762 8990 1764 9042
rect 1708 8372 1764 8990
rect 1932 8428 1988 19068
rect 2716 19012 2772 19022
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 2044 18228 2100 18510
rect 2492 18340 2548 18350
rect 2492 18246 2548 18284
rect 2044 18162 2100 18172
rect 2268 17668 2324 17678
rect 2268 17666 2436 17668
rect 2268 17614 2270 17666
rect 2322 17614 2436 17666
rect 2268 17612 2436 17614
rect 2268 17602 2324 17612
rect 2268 17444 2324 17454
rect 2268 16882 2324 17388
rect 2268 16830 2270 16882
rect 2322 16830 2324 16882
rect 2268 16818 2324 16830
rect 2380 16884 2436 17612
rect 2492 16884 2548 16894
rect 2380 16828 2492 16884
rect 2492 15314 2548 16828
rect 2492 15262 2494 15314
rect 2546 15262 2548 15314
rect 2492 15250 2548 15262
rect 2604 16324 2660 16334
rect 2268 14532 2324 14542
rect 2268 14530 2436 14532
rect 2268 14478 2270 14530
rect 2322 14478 2436 14530
rect 2268 14476 2436 14478
rect 2268 14466 2324 14476
rect 2268 14196 2324 14206
rect 2156 14140 2268 14196
rect 2044 9268 2100 9278
rect 2044 9174 2100 9212
rect 2156 8428 2212 14140
rect 2268 14130 2324 14140
rect 2268 13748 2324 13758
rect 2268 13654 2324 13692
rect 2268 12068 2324 12078
rect 2268 11974 2324 12012
rect 2380 11508 2436 14476
rect 2380 11442 2436 11452
rect 2268 10724 2324 10734
rect 2268 10630 2324 10668
rect 2492 8930 2548 8942
rect 2492 8878 2494 8930
rect 2546 8878 2548 8930
rect 1932 8372 2100 8428
rect 2156 8372 2324 8428
rect 1708 8306 1764 8316
rect 2044 7698 2100 8372
rect 2044 7646 2046 7698
rect 2098 7646 2100 7698
rect 2044 7634 2100 7646
rect 1708 7474 1764 7486
rect 1708 7422 1710 7474
rect 1762 7422 1764 7474
rect 1708 7364 1764 7422
rect 1708 6804 1764 7308
rect 1708 6738 1764 6748
rect 2268 6132 2324 8372
rect 2492 8372 2548 8878
rect 2492 8306 2548 8316
rect 2492 7364 2548 7374
rect 2492 7270 2548 7308
rect 1932 6076 2324 6132
rect 1820 5906 1876 5918
rect 1820 5854 1822 5906
rect 1874 5854 1876 5906
rect 1820 5236 1876 5854
rect 1820 5142 1876 5180
rect 1708 4338 1764 4350
rect 1708 4286 1710 4338
rect 1762 4286 1764 4338
rect 1708 4228 1764 4286
rect 1708 3668 1764 4172
rect 1708 3602 1764 3612
rect 1708 3442 1764 3454
rect 1708 3390 1710 3442
rect 1762 3390 1764 3442
rect 1708 3332 1764 3390
rect 1932 3444 1988 6076
rect 2268 5908 2324 5918
rect 2604 5908 2660 16268
rect 2268 5906 2660 5908
rect 2268 5854 2270 5906
rect 2322 5854 2660 5906
rect 2268 5852 2660 5854
rect 2268 5842 2324 5852
rect 2716 5684 2772 18956
rect 2940 17556 2996 17566
rect 2940 17462 2996 17500
rect 3052 10724 3108 34188
rect 3164 23268 3220 34972
rect 3276 34914 3332 35308
rect 3276 34862 3278 34914
rect 3330 34862 3332 34914
rect 3276 34580 3332 34862
rect 3500 34692 3556 35868
rect 3612 34916 3668 34954
rect 3612 34850 3668 34860
rect 3612 34692 3668 34702
rect 3500 34690 3668 34692
rect 3500 34638 3614 34690
rect 3666 34638 3668 34690
rect 3500 34636 3668 34638
rect 3612 34626 3668 34636
rect 3276 34524 3444 34580
rect 3388 34468 3444 34524
rect 3388 34412 3668 34468
rect 3388 34020 3444 34030
rect 3612 34020 3668 34412
rect 3388 34018 3556 34020
rect 3388 33966 3390 34018
rect 3442 33966 3556 34018
rect 3388 33964 3556 33966
rect 3388 33954 3444 33964
rect 3164 23202 3220 23212
rect 3500 33796 3556 33964
rect 3612 33954 3668 33964
rect 3724 34018 3780 37998
rect 3836 38050 3892 38220
rect 3836 37998 3838 38050
rect 3890 37998 3892 38050
rect 3836 37986 3892 37998
rect 4060 36596 4116 44158
rect 4284 44100 4340 44110
rect 4284 43538 4340 44044
rect 4284 43486 4286 43538
rect 4338 43486 4340 43538
rect 4284 43474 4340 43486
rect 4732 43540 4788 44380
rect 4844 44324 4900 44334
rect 4844 44230 4900 44268
rect 4956 43988 5012 45614
rect 4956 43922 5012 43932
rect 5292 43764 5348 43774
rect 5404 43764 5460 45836
rect 5628 46900 5684 46910
rect 5628 46004 5684 46844
rect 6748 46788 6804 49200
rect 6748 46732 7252 46788
rect 5628 45890 5684 45948
rect 6636 46004 6692 46014
rect 6636 45910 6692 45948
rect 7196 46004 7252 46732
rect 7196 46002 7588 46004
rect 7196 45950 7198 46002
rect 7250 45950 7588 46002
rect 7196 45948 7588 45950
rect 7196 45938 7252 45948
rect 5628 45838 5630 45890
rect 5682 45838 5684 45890
rect 5628 45826 5684 45838
rect 6188 45890 6244 45902
rect 6188 45838 6190 45890
rect 6242 45838 6244 45890
rect 5292 43762 5460 43764
rect 5292 43710 5294 43762
rect 5346 43710 5460 43762
rect 5292 43708 5460 43710
rect 5628 44324 5684 44334
rect 5628 43764 5684 44268
rect 5964 44324 6020 44334
rect 5964 44230 6020 44268
rect 5292 43698 5348 43708
rect 4732 43538 4900 43540
rect 4732 43486 4734 43538
rect 4786 43486 4900 43538
rect 4732 43484 4900 43486
rect 4732 43446 4788 43484
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4284 42756 4340 42766
rect 4284 42662 4340 42700
rect 4732 42756 4788 42766
rect 4844 42756 4900 43484
rect 4732 42754 4900 42756
rect 4732 42702 4734 42754
rect 4786 42702 4900 42754
rect 4732 42700 4900 42702
rect 5628 43426 5684 43708
rect 5628 43374 5630 43426
rect 5682 43374 5684 43426
rect 4732 42690 4788 42700
rect 4956 42530 5012 42542
rect 4956 42478 4958 42530
rect 5010 42478 5012 42530
rect 4508 41860 4564 41870
rect 4508 41766 4564 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4844 41300 4900 41310
rect 4844 41206 4900 41244
rect 4284 40402 4340 40414
rect 4284 40350 4286 40402
rect 4338 40350 4340 40402
rect 4284 40292 4340 40350
rect 4284 40226 4340 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4284 38834 4340 38846
rect 4284 38782 4286 38834
rect 4338 38782 4340 38834
rect 4284 38052 4340 38782
rect 4844 38724 4900 38734
rect 4844 38630 4900 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4956 38164 5012 42478
rect 5516 41300 5572 41310
rect 5292 39508 5348 39518
rect 5180 38724 5236 38734
rect 4956 38098 5012 38108
rect 5068 38722 5236 38724
rect 5068 38670 5182 38722
rect 5234 38670 5236 38722
rect 5068 38668 5236 38670
rect 4284 37986 4340 37996
rect 4508 37938 4564 37950
rect 4844 37940 4900 37950
rect 4508 37886 4510 37938
rect 4562 37886 4564 37938
rect 4396 37828 4452 37838
rect 4060 36530 4116 36540
rect 4172 37826 4452 37828
rect 4172 37774 4398 37826
rect 4450 37774 4452 37826
rect 4172 37772 4452 37774
rect 4172 36260 4228 37772
rect 4396 37762 4452 37772
rect 4284 37156 4340 37166
rect 4284 36482 4340 37100
rect 4508 37044 4564 37886
rect 4732 37884 4844 37940
rect 4732 37044 4788 37884
rect 4844 37846 4900 37884
rect 4956 37828 5012 37838
rect 5068 37828 5124 38668
rect 5180 38658 5236 38668
rect 5180 38052 5236 38062
rect 5292 38052 5348 39452
rect 5180 38050 5348 38052
rect 5180 37998 5182 38050
rect 5234 37998 5348 38050
rect 5180 37996 5348 37998
rect 5180 37986 5236 37996
rect 4956 37826 5124 37828
rect 4956 37774 4958 37826
rect 5010 37774 5124 37826
rect 4956 37772 5124 37774
rect 4956 37762 5012 37772
rect 4844 37604 4900 37614
rect 4900 37548 5012 37604
rect 4844 37538 4900 37548
rect 4732 36988 4900 37044
rect 4508 36978 4564 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 36820 4900 36988
rect 4844 36596 4900 36764
rect 4956 36706 5012 37548
rect 5068 37492 5124 37772
rect 5180 37492 5236 37502
rect 5068 37436 5180 37492
rect 5180 37426 5236 37436
rect 5180 37154 5236 37166
rect 5180 37102 5182 37154
rect 5234 37102 5236 37154
rect 5180 37044 5236 37102
rect 5180 36978 5236 36988
rect 4956 36654 4958 36706
rect 5010 36654 5012 36706
rect 4956 36642 5012 36654
rect 4284 36430 4286 36482
rect 4338 36430 4340 36482
rect 4284 36418 4340 36430
rect 4620 36540 4900 36596
rect 3836 36204 4228 36260
rect 3836 34914 3892 36204
rect 4620 35924 4676 36540
rect 4956 36484 5012 36494
rect 3836 34862 3838 34914
rect 3890 34862 3892 34914
rect 3836 34850 3892 34862
rect 4060 35922 4676 35924
rect 4060 35870 4622 35922
rect 4674 35870 4676 35922
rect 4060 35868 4676 35870
rect 4060 34914 4116 35868
rect 4620 35858 4676 35868
rect 4844 36428 4956 36484
rect 4284 35698 4340 35710
rect 4284 35646 4286 35698
rect 4338 35646 4340 35698
rect 4284 35140 4340 35646
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4284 35074 4340 35084
rect 4732 35140 4788 35150
rect 4844 35140 4900 36428
rect 4956 36418 5012 36428
rect 5068 36372 5124 36382
rect 5068 36278 5124 36316
rect 5516 36372 5572 41244
rect 5628 40964 5684 43374
rect 5740 40964 5796 40974
rect 5684 40962 5796 40964
rect 5684 40910 5742 40962
rect 5794 40910 5796 40962
rect 5684 40908 5796 40910
rect 5628 37268 5684 40908
rect 5740 40898 5796 40908
rect 5628 37174 5684 37212
rect 5628 36820 5684 36830
rect 5628 36482 5684 36764
rect 5852 36708 5908 36718
rect 5740 36596 5796 36606
rect 5740 36502 5796 36540
rect 5628 36430 5630 36482
rect 5682 36430 5684 36482
rect 5628 36418 5684 36430
rect 5852 36482 5908 36652
rect 5852 36430 5854 36482
rect 5906 36430 5908 36482
rect 5852 36418 5908 36430
rect 6076 36484 6132 36494
rect 6076 36390 6132 36428
rect 5516 36306 5572 36316
rect 6188 35812 6244 45838
rect 7196 45668 7252 45678
rect 7196 45106 7252 45612
rect 7532 45218 7588 45948
rect 8092 46002 8148 49200
rect 8092 45950 8094 46002
rect 8146 45950 8148 46002
rect 8092 45444 8148 45950
rect 9436 45892 9492 49200
rect 10780 46004 10836 49200
rect 10780 46002 11060 46004
rect 10780 45950 10782 46002
rect 10834 45950 11060 46002
rect 10780 45948 11060 45950
rect 10780 45938 10836 45948
rect 9660 45892 9716 45902
rect 9436 45890 9716 45892
rect 9436 45838 9662 45890
rect 9714 45838 9716 45890
rect 9436 45836 9716 45838
rect 8764 45778 8820 45790
rect 8764 45726 8766 45778
rect 8818 45726 8820 45778
rect 8428 45668 8484 45678
rect 8428 45574 8484 45612
rect 8092 45388 8484 45444
rect 7532 45166 7534 45218
rect 7586 45166 7588 45218
rect 7532 45154 7588 45166
rect 7868 45220 7924 45230
rect 7868 45126 7924 45164
rect 7196 45054 7198 45106
rect 7250 45054 7252 45106
rect 7196 45042 7252 45054
rect 8428 45106 8484 45388
rect 8652 45220 8708 45230
rect 8652 45126 8708 45164
rect 8428 45054 8430 45106
rect 8482 45054 8484 45106
rect 8428 45042 8484 45054
rect 8092 44436 8148 44446
rect 8764 44436 8820 45726
rect 9660 45330 9716 45836
rect 11004 45890 11060 45948
rect 11004 45838 11006 45890
rect 11058 45838 11060 45890
rect 11004 45826 11060 45838
rect 12124 45892 12180 49200
rect 13468 46004 13524 49200
rect 14812 46004 14868 49200
rect 16156 46004 16212 49200
rect 16380 46004 16436 46014
rect 13468 46002 13748 46004
rect 13468 45950 13470 46002
rect 13522 45950 13748 46002
rect 13468 45948 13748 45950
rect 13468 45938 13524 45948
rect 12236 45892 12292 45902
rect 12124 45890 12852 45892
rect 12124 45838 12238 45890
rect 12290 45838 12852 45890
rect 12124 45836 12852 45838
rect 12236 45826 12292 45836
rect 9996 45668 10052 45678
rect 11340 45668 11396 45678
rect 9660 45278 9662 45330
rect 9714 45278 9716 45330
rect 9660 45266 9716 45278
rect 9772 45666 10052 45668
rect 9772 45614 9998 45666
rect 10050 45614 10052 45666
rect 9772 45612 10052 45614
rect 8876 44436 8932 44446
rect 8764 44434 8932 44436
rect 8764 44382 8878 44434
rect 8930 44382 8932 44434
rect 8764 44380 8932 44382
rect 6748 44212 6804 44222
rect 6748 44210 8036 44212
rect 6748 44158 6750 44210
rect 6802 44158 8036 44210
rect 6748 44156 8036 44158
rect 6748 44146 6804 44156
rect 7420 43988 7476 43998
rect 6748 43650 6804 43662
rect 6748 43598 6750 43650
rect 6802 43598 6804 43650
rect 6748 42756 6804 43598
rect 7420 43650 7476 43932
rect 7420 43598 7422 43650
rect 7474 43598 7476 43650
rect 7420 43586 7476 43598
rect 6748 42690 6804 42700
rect 6972 43538 7028 43550
rect 6972 43486 6974 43538
rect 7026 43486 7028 43538
rect 6636 41858 6692 41870
rect 6636 41806 6638 41858
rect 6690 41806 6692 41858
rect 6636 40516 6692 41806
rect 6972 41300 7028 43486
rect 7868 43538 7924 43550
rect 7868 43486 7870 43538
rect 7922 43486 7924 43538
rect 7532 43314 7588 43326
rect 7532 43262 7534 43314
rect 7586 43262 7588 43314
rect 7084 41972 7140 41982
rect 7308 41972 7364 41982
rect 7084 41970 7252 41972
rect 7084 41918 7086 41970
rect 7138 41918 7252 41970
rect 7084 41916 7252 41918
rect 7084 41906 7140 41916
rect 6972 41234 7028 41244
rect 6860 40964 6916 40974
rect 6860 40870 6916 40908
rect 6636 40450 6692 40460
rect 6748 40514 6804 40526
rect 6748 40462 6750 40514
rect 6802 40462 6804 40514
rect 6748 40292 6804 40462
rect 7084 40516 7140 40526
rect 7196 40516 7252 41916
rect 7308 41878 7364 41916
rect 7420 41860 7476 41870
rect 7420 41766 7476 41804
rect 7196 40460 7364 40516
rect 7084 40422 7140 40460
rect 6748 40226 6804 40236
rect 7196 39956 7252 39966
rect 7084 39620 7140 39630
rect 7196 39620 7252 39900
rect 7084 39618 7252 39620
rect 7084 39566 7086 39618
rect 7138 39566 7252 39618
rect 7084 39564 7252 39566
rect 7308 39620 7364 40460
rect 7084 39554 7140 39564
rect 7308 39526 7364 39564
rect 6748 39508 6804 39518
rect 6748 39414 6804 39452
rect 6972 39394 7028 39406
rect 6972 39342 6974 39394
rect 7026 39342 7028 39394
rect 6972 39060 7028 39342
rect 6972 39004 7364 39060
rect 7308 38946 7364 39004
rect 7308 38894 7310 38946
rect 7362 38894 7364 38946
rect 7308 38882 7364 38894
rect 6412 36482 6468 36494
rect 6412 36430 6414 36482
rect 6466 36430 6468 36482
rect 6412 36260 6468 36430
rect 6860 36260 6916 36270
rect 6412 36258 6916 36260
rect 6412 36206 6862 36258
rect 6914 36206 6916 36258
rect 6412 36204 6916 36206
rect 6188 35746 6244 35756
rect 4732 35138 4900 35140
rect 4732 35086 4734 35138
rect 4786 35086 4900 35138
rect 4732 35084 4900 35086
rect 4956 35698 5012 35710
rect 4956 35646 4958 35698
rect 5010 35646 5012 35698
rect 4732 35074 4788 35084
rect 4060 34862 4062 34914
rect 4114 34862 4116 34914
rect 4060 34850 4116 34862
rect 4396 34804 4452 34814
rect 4172 34748 4396 34804
rect 3724 33966 3726 34018
rect 3778 33966 3780 34018
rect 3724 33954 3780 33966
rect 3836 34242 3892 34254
rect 3836 34190 3838 34242
rect 3890 34190 3892 34242
rect 3836 33796 3892 34190
rect 4060 34244 4116 34254
rect 4172 34244 4228 34748
rect 4396 34710 4452 34748
rect 4844 34804 4900 34814
rect 4956 34804 5012 35646
rect 6636 35028 6692 35038
rect 4900 34748 5012 34804
rect 5628 34804 5684 34814
rect 4844 34738 4900 34748
rect 5628 34710 5684 34748
rect 5964 34804 6020 34814
rect 5964 34710 6020 34748
rect 4060 34242 4228 34244
rect 4060 34190 4062 34242
rect 4114 34190 4228 34242
rect 4060 34188 4228 34190
rect 4620 34690 4676 34702
rect 4620 34638 4622 34690
rect 4674 34638 4676 34690
rect 4060 34178 4116 34188
rect 4508 34020 4564 34030
rect 4508 33926 4564 33964
rect 4284 33908 4340 33918
rect 3500 33740 3892 33796
rect 4172 33906 4340 33908
rect 4172 33854 4286 33906
rect 4338 33854 4340 33906
rect 4172 33852 4340 33854
rect 3388 16884 3444 16894
rect 3388 16790 3444 16828
rect 3500 16548 3556 33740
rect 4060 31668 4116 31678
rect 4060 31574 4116 31612
rect 4172 31444 4228 33852
rect 4284 33842 4340 33852
rect 4620 33906 4676 34638
rect 4620 33854 4622 33906
rect 4674 33854 4676 33906
rect 4620 33842 4676 33854
rect 4956 34018 5012 34030
rect 4956 33966 4958 34018
rect 5010 33966 5012 34018
rect 4956 33906 5012 33966
rect 4956 33854 4958 33906
rect 5010 33854 5012 33906
rect 4956 33842 5012 33854
rect 6412 33796 6468 33806
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 32562 4340 32574
rect 4284 32510 4286 32562
rect 4338 32510 4340 32562
rect 4284 31780 4340 32510
rect 5068 32450 5124 32462
rect 5068 32398 5070 32450
rect 5122 32398 5124 32450
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5068 31892 5124 32398
rect 4284 31714 4340 31724
rect 4844 31836 5068 31892
rect 4844 31778 4900 31836
rect 4844 31726 4846 31778
rect 4898 31726 4900 31778
rect 4844 31714 4900 31726
rect 4060 31388 4228 31444
rect 3948 30884 4004 30894
rect 3948 30210 4004 30828
rect 3948 30158 3950 30210
rect 4002 30158 4004 30210
rect 3948 30146 4004 30158
rect 4060 28420 4116 31388
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 29426 4340 29438
rect 4284 29374 4286 29426
rect 4338 29374 4340 29426
rect 4172 28868 4228 28878
rect 4172 28532 4228 28812
rect 4284 28756 4340 29374
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4284 28690 4340 28700
rect 5068 28756 5124 31836
rect 5740 31780 5796 31790
rect 5740 31686 5796 31724
rect 5852 31556 5908 31566
rect 5852 31462 5908 31500
rect 6076 31220 6132 31230
rect 6076 31106 6132 31164
rect 6076 31054 6078 31106
rect 6130 31054 6132 31106
rect 6076 31042 6132 31054
rect 5740 28756 5796 28766
rect 5068 28754 5796 28756
rect 5068 28702 5742 28754
rect 5794 28702 5796 28754
rect 5068 28700 5796 28702
rect 5068 28642 5124 28700
rect 5068 28590 5070 28642
rect 5122 28590 5124 28642
rect 5068 28578 5124 28590
rect 4284 28532 4340 28542
rect 4172 28530 4340 28532
rect 4172 28478 4286 28530
rect 4338 28478 4340 28530
rect 4172 28476 4340 28478
rect 4284 28466 4340 28476
rect 4060 28364 4228 28420
rect 4060 27860 4116 27870
rect 4060 26290 4116 27804
rect 4060 26238 4062 26290
rect 4114 26238 4116 26290
rect 4060 26226 4116 26238
rect 4172 26068 4228 28364
rect 5068 28084 5124 28094
rect 5068 27970 5124 28028
rect 5068 27918 5070 27970
rect 5122 27918 5124 27970
rect 5068 27906 5124 27918
rect 4284 27636 4340 27646
rect 4284 27186 4340 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27134 4286 27186
rect 4338 27134 4340 27186
rect 4284 27122 4340 27134
rect 5068 27076 5124 27086
rect 5180 27076 5236 28700
rect 5740 28084 5796 28700
rect 6300 28084 6356 28094
rect 5740 28082 6356 28084
rect 5740 28030 6302 28082
rect 6354 28030 6356 28082
rect 5740 28028 6356 28030
rect 5740 27858 5796 28028
rect 5740 27806 5742 27858
rect 5794 27806 5796 27858
rect 5740 27794 5796 27806
rect 5852 27186 5908 28028
rect 6300 28018 6356 28028
rect 5852 27134 5854 27186
rect 5906 27134 5908 27186
rect 5852 27122 5908 27134
rect 5068 27074 5236 27076
rect 5068 27022 5070 27074
rect 5122 27022 5236 27074
rect 5068 27020 5236 27022
rect 5068 27010 5124 27020
rect 4508 26964 4564 26974
rect 3948 26012 4228 26068
rect 4284 26852 4564 26908
rect 3948 17220 4004 26012
rect 4284 25506 4340 26852
rect 4956 26180 5012 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 25442 4340 25454
rect 4956 24834 5012 26124
rect 6412 24948 6468 33740
rect 6636 31892 6692 34972
rect 6860 33236 6916 36204
rect 7308 35364 7364 35374
rect 7196 35308 7308 35364
rect 7196 34804 7252 35308
rect 7308 35298 7364 35308
rect 7308 35140 7364 35150
rect 7308 35046 7364 35084
rect 7308 34804 7364 34814
rect 7196 34802 7364 34804
rect 7196 34750 7310 34802
rect 7362 34750 7364 34802
rect 7196 34748 7364 34750
rect 7308 34738 7364 34748
rect 7420 34802 7476 34814
rect 7420 34750 7422 34802
rect 7474 34750 7476 34802
rect 7420 34692 7476 34750
rect 7532 34692 7588 43262
rect 7756 42644 7812 42654
rect 7756 42550 7812 42588
rect 7644 42532 7700 42542
rect 7644 41970 7700 42476
rect 7868 42082 7924 43486
rect 7868 42030 7870 42082
rect 7922 42030 7924 42082
rect 7868 42018 7924 42030
rect 7644 41918 7646 41970
rect 7698 41918 7700 41970
rect 7644 41906 7700 41918
rect 7980 41970 8036 44156
rect 8092 43988 8148 44380
rect 8092 43922 8148 43932
rect 8876 43708 8932 44380
rect 9324 44098 9380 44110
rect 9324 44046 9326 44098
rect 9378 44046 9380 44098
rect 9324 43708 9380 44046
rect 8092 43650 8148 43662
rect 8876 43652 9044 43708
rect 8092 43598 8094 43650
rect 8146 43598 8148 43650
rect 8092 42868 8148 43598
rect 8092 42802 8148 42812
rect 8204 43538 8260 43550
rect 8204 43486 8206 43538
rect 8258 43486 8260 43538
rect 8092 42644 8148 42682
rect 8092 42578 8148 42588
rect 7980 41918 7982 41970
rect 8034 41918 8036 41970
rect 7980 41906 8036 41918
rect 8092 42420 8148 42430
rect 8204 42420 8260 43486
rect 8988 42868 9044 43652
rect 9324 43652 9604 43708
rect 9324 43586 9380 43596
rect 8764 42756 8820 42766
rect 8764 42662 8820 42700
rect 8428 42532 8484 42542
rect 8652 42532 8708 42542
rect 8428 42438 8484 42476
rect 8540 42530 8708 42532
rect 8540 42478 8654 42530
rect 8706 42478 8708 42530
rect 8540 42476 8708 42478
rect 8148 42364 8260 42420
rect 8092 41074 8148 42364
rect 8428 42084 8484 42094
rect 8428 41990 8484 42028
rect 8204 41970 8260 41982
rect 8204 41918 8206 41970
rect 8258 41918 8260 41970
rect 8204 41860 8260 41918
rect 8540 41860 8596 42476
rect 8652 42466 8708 42476
rect 8988 42532 9044 42812
rect 9436 43428 9492 43438
rect 8988 42466 9044 42476
rect 9324 42530 9380 42542
rect 9324 42478 9326 42530
rect 9378 42478 9380 42530
rect 8876 42082 8932 42094
rect 8876 42030 8878 42082
rect 8930 42030 8932 42082
rect 8652 41972 8708 41982
rect 8652 41878 8708 41916
rect 8204 41794 8260 41804
rect 8428 41804 8596 41860
rect 8092 41022 8094 41074
rect 8146 41022 8148 41074
rect 8092 41010 8148 41022
rect 8316 41186 8372 41198
rect 8316 41134 8318 41186
rect 8370 41134 8372 41186
rect 8204 40402 8260 40414
rect 8204 40350 8206 40402
rect 8258 40350 8260 40402
rect 8204 39956 8260 40350
rect 8204 39890 8260 39900
rect 8316 39172 8372 41134
rect 8428 40740 8484 41804
rect 8876 41300 8932 42030
rect 9324 42084 9380 42478
rect 8876 41234 8932 41244
rect 8988 41970 9044 41982
rect 8988 41918 8990 41970
rect 9042 41918 9044 41970
rect 8988 41188 9044 41918
rect 9212 41300 9268 41310
rect 9212 41206 9268 41244
rect 8988 41076 9044 41132
rect 8428 40674 8484 40684
rect 8540 41020 9044 41076
rect 8428 40514 8484 40526
rect 8428 40462 8430 40514
rect 8482 40462 8484 40514
rect 8428 40404 8484 40462
rect 8540 40514 8596 41020
rect 8540 40462 8542 40514
rect 8594 40462 8596 40514
rect 8540 40450 8596 40462
rect 8988 40740 9044 40750
rect 8988 40626 9044 40684
rect 8988 40574 8990 40626
rect 9042 40574 9044 40626
rect 8428 40338 8484 40348
rect 8988 40404 9044 40574
rect 8988 40338 9044 40348
rect 7980 39116 8372 39172
rect 7980 38668 8036 39116
rect 8540 39060 8596 39070
rect 8092 39004 8540 39060
rect 8092 38834 8148 39004
rect 8092 38782 8094 38834
rect 8146 38782 8148 38834
rect 8092 38770 8148 38782
rect 7868 38612 8036 38668
rect 8540 38722 8596 39004
rect 8540 38670 8542 38722
rect 8594 38670 8596 38722
rect 7644 38052 7700 38062
rect 7644 37490 7700 37996
rect 7644 37438 7646 37490
rect 7698 37438 7700 37490
rect 7644 37426 7700 37438
rect 7756 37826 7812 37838
rect 7756 37774 7758 37826
rect 7810 37774 7812 37826
rect 7756 37156 7812 37774
rect 7756 37090 7812 37100
rect 7868 36932 7924 38612
rect 8092 37938 8148 37950
rect 8092 37886 8094 37938
rect 8146 37886 8148 37938
rect 8092 37492 8148 37886
rect 8092 37426 8148 37436
rect 7980 37268 8036 37278
rect 7980 37266 8148 37268
rect 7980 37214 7982 37266
rect 8034 37214 8148 37266
rect 7980 37212 8148 37214
rect 7980 37202 8036 37212
rect 8092 37044 8148 37212
rect 8092 36978 8148 36988
rect 7868 36876 8036 36932
rect 7980 34804 8036 36876
rect 8316 36484 8372 36494
rect 7868 34692 7924 34702
rect 7420 34690 7924 34692
rect 7420 34638 7870 34690
rect 7922 34638 7924 34690
rect 7420 34636 7924 34638
rect 7420 33796 7476 34636
rect 7868 34626 7924 34636
rect 7420 33730 7476 33740
rect 7644 34020 7700 34030
rect 6860 33180 7476 33236
rect 6636 30996 6692 31836
rect 6748 30996 6804 31006
rect 7308 30996 7364 31006
rect 6636 30994 7364 30996
rect 6636 30942 6750 30994
rect 6802 30942 7310 30994
rect 7362 30942 7364 30994
rect 6636 30940 7364 30942
rect 6748 30930 6804 30940
rect 7308 30930 7364 30940
rect 6412 24882 6468 24892
rect 6524 30436 6580 30446
rect 4956 24782 4958 24834
rect 5010 24782 5012 24834
rect 4956 24770 5012 24782
rect 5740 24722 5796 24734
rect 5740 24670 5742 24722
rect 5794 24670 5796 24722
rect 4284 24612 4340 24622
rect 5740 24612 5796 24670
rect 6300 24612 6356 24622
rect 5740 24610 6356 24612
rect 5740 24558 6302 24610
rect 6354 24558 6356 24610
rect 5740 24556 6356 24558
rect 4284 23940 4340 24556
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23846 4340 23884
rect 5964 23604 6020 23614
rect 4284 23268 4340 23278
rect 4284 23154 4340 23212
rect 5740 23268 5796 23278
rect 5740 23174 5796 23212
rect 4284 23102 4286 23154
rect 4338 23102 4340 23154
rect 4284 23090 4340 23102
rect 5852 23156 5908 23166
rect 5852 23062 5908 23100
rect 5180 23044 5236 23054
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4508 22596 4564 22606
rect 4172 22484 4228 22494
rect 4172 22390 4228 22428
rect 4396 21588 4452 21598
rect 4508 21588 4564 22540
rect 4956 22372 5012 22382
rect 5180 22372 5236 22988
rect 5964 22594 6020 23548
rect 6300 23044 6356 24556
rect 6524 23548 6580 30380
rect 6860 27300 6916 27310
rect 6860 27206 6916 27244
rect 6748 26964 6804 27002
rect 6748 26898 6804 26908
rect 7420 26852 7476 33180
rect 7644 31444 7700 33964
rect 7980 33348 8036 34748
rect 7980 33282 8036 33292
rect 8204 36370 8260 36382
rect 8204 36318 8206 36370
rect 8258 36318 8260 36370
rect 8204 32004 8260 36318
rect 8316 35364 8372 36428
rect 8428 36372 8484 36382
rect 8428 36278 8484 36316
rect 8316 35026 8372 35308
rect 8316 34974 8318 35026
rect 8370 34974 8372 35026
rect 8316 34962 8372 34974
rect 8540 35028 8596 38670
rect 8876 37156 8932 37166
rect 8876 36482 8932 37100
rect 8876 36430 8878 36482
rect 8930 36430 8932 36482
rect 8876 36418 8932 36430
rect 8540 34962 8596 34972
rect 8652 36258 8708 36270
rect 8652 36206 8654 36258
rect 8706 36206 8708 36258
rect 8652 34916 8708 36206
rect 9324 35924 9380 42028
rect 9436 39060 9492 43372
rect 9548 42644 9604 43652
rect 9548 42578 9604 42588
rect 9436 38994 9492 39004
rect 9660 42532 9716 42542
rect 9212 35868 9380 35924
rect 9436 37490 9492 37502
rect 9436 37438 9438 37490
rect 9490 37438 9492 37490
rect 8988 34916 9044 34926
rect 8652 34914 9044 34916
rect 8652 34862 8990 34914
rect 9042 34862 9044 34914
rect 8652 34860 9044 34862
rect 8988 34850 9044 34860
rect 8204 31938 8260 31948
rect 8764 34690 8820 34702
rect 8764 34638 8766 34690
rect 8818 34638 8820 34690
rect 7644 31378 7700 31388
rect 7980 31668 8036 31678
rect 7980 31218 8036 31612
rect 7980 31166 7982 31218
rect 8034 31166 8036 31218
rect 7980 31154 8036 31166
rect 8092 31556 8148 31566
rect 8092 31106 8148 31500
rect 8316 31556 8372 31566
rect 8316 31462 8372 31500
rect 8540 31556 8596 31566
rect 8540 31462 8596 31500
rect 8764 31332 8820 34638
rect 9212 32340 9268 35868
rect 9436 35028 9492 37438
rect 9548 37380 9604 37418
rect 9548 37314 9604 37324
rect 9548 37156 9604 37166
rect 9548 36482 9604 37100
rect 9548 36430 9550 36482
rect 9602 36430 9604 36482
rect 9548 35922 9604 36430
rect 9660 36484 9716 42476
rect 9772 37156 9828 45612
rect 9996 45602 10052 45612
rect 11228 45666 11396 45668
rect 11228 45614 11342 45666
rect 11394 45614 11396 45666
rect 11228 45612 11396 45614
rect 10556 43652 10612 43662
rect 10556 43558 10612 43596
rect 10444 43540 10500 43550
rect 9996 43538 10500 43540
rect 9996 43486 10446 43538
rect 10498 43486 10500 43538
rect 9996 43484 10500 43486
rect 9884 42754 9940 42766
rect 9884 42702 9886 42754
rect 9938 42702 9940 42754
rect 9884 42644 9940 42702
rect 9884 42578 9940 42588
rect 9996 42756 10052 43484
rect 10444 43474 10500 43484
rect 10556 43316 10612 43326
rect 10556 43314 10724 43316
rect 10556 43262 10558 43314
rect 10610 43262 10724 43314
rect 10556 43260 10724 43262
rect 10556 43250 10612 43260
rect 9996 42420 10052 42700
rect 9884 42364 10052 42420
rect 10556 42642 10612 42654
rect 10556 42590 10558 42642
rect 10610 42590 10612 42642
rect 9884 42082 9940 42364
rect 10556 42194 10612 42590
rect 10556 42142 10558 42194
rect 10610 42142 10612 42194
rect 10556 42130 10612 42142
rect 9884 42030 9886 42082
rect 9938 42030 9940 42082
rect 9884 42018 9940 42030
rect 9996 42084 10052 42094
rect 9996 41990 10052 42028
rect 10220 42082 10276 42094
rect 10220 42030 10222 42082
rect 10274 42030 10276 42082
rect 10220 41972 10276 42030
rect 10332 41972 10388 41982
rect 10220 41970 10388 41972
rect 10220 41918 10334 41970
rect 10386 41918 10388 41970
rect 10220 41916 10388 41918
rect 10332 41906 10388 41916
rect 10668 41972 10724 43260
rect 11116 43092 11172 43102
rect 11004 43036 11116 43092
rect 10668 41906 10724 41916
rect 10780 41970 10836 41982
rect 10780 41918 10782 41970
rect 10834 41918 10836 41970
rect 10780 41412 10836 41918
rect 10780 41346 10836 41356
rect 10892 41970 10948 41982
rect 10892 41918 10894 41970
rect 10946 41918 10948 41970
rect 10892 41748 10948 41918
rect 10668 40516 10724 40526
rect 10220 39620 10276 39630
rect 10220 39058 10276 39564
rect 10220 39006 10222 39058
rect 10274 39006 10276 39058
rect 10220 38994 10276 39006
rect 9884 38836 9940 38846
rect 9884 38742 9940 38780
rect 10556 38836 10612 38846
rect 10556 38742 10612 38780
rect 9996 38276 10052 38286
rect 9996 38050 10052 38220
rect 9996 37998 9998 38050
rect 10050 37998 10052 38050
rect 9996 37986 10052 37998
rect 10444 38164 10500 38174
rect 10444 38050 10500 38108
rect 10444 37998 10446 38050
rect 10498 37998 10500 38050
rect 10444 37986 10500 37998
rect 10220 37826 10276 37838
rect 10220 37774 10222 37826
rect 10274 37774 10276 37826
rect 9996 37380 10052 37390
rect 9772 37090 9828 37100
rect 9884 37266 9940 37278
rect 9884 37214 9886 37266
rect 9938 37214 9940 37266
rect 9772 36484 9828 36494
rect 9660 36482 9828 36484
rect 9660 36430 9774 36482
rect 9826 36430 9828 36482
rect 9660 36428 9828 36430
rect 9772 36418 9828 36428
rect 9884 36484 9940 37214
rect 9884 36418 9940 36428
rect 9996 36482 10052 37324
rect 10220 37268 10276 37774
rect 10220 37202 10276 37212
rect 10332 37826 10388 37838
rect 10332 37774 10334 37826
rect 10386 37774 10388 37826
rect 9996 36430 9998 36482
rect 10050 36430 10052 36482
rect 9996 36418 10052 36430
rect 10220 36370 10276 36382
rect 10220 36318 10222 36370
rect 10274 36318 10276 36370
rect 9884 36260 9940 36270
rect 9548 35870 9550 35922
rect 9602 35870 9604 35922
rect 9548 35858 9604 35870
rect 9660 36258 9940 36260
rect 9660 36206 9886 36258
rect 9938 36206 9940 36258
rect 9660 36204 9940 36206
rect 9660 35476 9716 36204
rect 9884 36194 9940 36204
rect 9212 32274 9268 32284
rect 9324 34972 9492 35028
rect 9548 35420 9716 35476
rect 9884 35700 9940 35710
rect 9324 32116 9380 34972
rect 9436 34804 9492 34814
rect 9436 34710 9492 34748
rect 9548 33572 9604 35420
rect 9884 35308 9940 35644
rect 10220 35588 10276 36318
rect 10332 35924 10388 37774
rect 10556 37826 10612 37838
rect 10556 37774 10558 37826
rect 10610 37774 10612 37826
rect 10556 36932 10612 37774
rect 10668 37266 10724 40460
rect 10892 39620 10948 41692
rect 10892 39554 10948 39564
rect 11004 38668 11060 43036
rect 11116 43026 11172 43036
rect 10668 37214 10670 37266
rect 10722 37214 10724 37266
rect 10668 37202 10724 37214
rect 10780 38612 11060 38668
rect 10668 36932 10724 36942
rect 10556 36876 10668 36932
rect 10668 36866 10724 36876
rect 10332 35858 10388 35868
rect 10668 36258 10724 36270
rect 10668 36206 10670 36258
rect 10722 36206 10724 36258
rect 10668 35700 10724 36206
rect 10668 35634 10724 35644
rect 10444 35588 10500 35598
rect 10220 35586 10500 35588
rect 10220 35534 10446 35586
rect 10498 35534 10500 35586
rect 10220 35532 10500 35534
rect 9660 35252 9716 35262
rect 9884 35252 10164 35308
rect 9660 34802 9716 35196
rect 9772 35140 9828 35150
rect 9772 34914 9828 35084
rect 9772 34862 9774 34914
rect 9826 34862 9828 34914
rect 9772 34850 9828 34862
rect 9660 34750 9662 34802
rect 9714 34750 9716 34802
rect 9660 34738 9716 34750
rect 9436 33516 9604 33572
rect 9436 33012 9492 33516
rect 9548 33348 9604 33358
rect 9548 33254 9604 33292
rect 9772 33348 9828 33358
rect 9772 33234 9828 33292
rect 10108 33348 10164 35252
rect 10444 34356 10500 35532
rect 10108 33282 10164 33292
rect 10220 34300 10500 34356
rect 9772 33182 9774 33234
rect 9826 33182 9828 33234
rect 9772 33170 9828 33182
rect 9884 33234 9940 33246
rect 9884 33182 9886 33234
rect 9938 33182 9940 33234
rect 9884 33124 9940 33182
rect 9884 33058 9940 33068
rect 9436 32956 9604 33012
rect 9100 32060 9380 32116
rect 9100 31890 9156 32060
rect 9436 32004 9492 32014
rect 9100 31838 9102 31890
rect 9154 31838 9156 31890
rect 9100 31826 9156 31838
rect 9212 31948 9436 32004
rect 8876 31778 8932 31790
rect 8876 31726 8878 31778
rect 8930 31726 8932 31778
rect 8876 31556 8932 31726
rect 8876 31490 8932 31500
rect 8764 31266 8820 31276
rect 8092 31054 8094 31106
rect 8146 31054 8148 31106
rect 8092 31042 8148 31054
rect 9100 31108 9156 31118
rect 7756 30996 7812 31006
rect 7756 30902 7812 30940
rect 8764 30996 8820 31006
rect 8764 30994 8932 30996
rect 8764 30942 8766 30994
rect 8818 30942 8932 30994
rect 8764 30940 8932 30942
rect 8764 30930 8820 30940
rect 7644 30884 7700 30894
rect 7644 30790 7700 30828
rect 8316 30882 8372 30894
rect 8316 30830 8318 30882
rect 8370 30830 8372 30882
rect 7980 30324 8036 30334
rect 7532 28756 7588 28766
rect 7532 28662 7588 28700
rect 7644 28644 7700 28654
rect 7644 28550 7700 28588
rect 7644 27860 7700 27870
rect 7644 27746 7700 27804
rect 7644 27694 7646 27746
rect 7698 27694 7700 27746
rect 7644 27682 7700 27694
rect 7756 27748 7812 27758
rect 7756 27654 7812 27692
rect 7420 26786 7476 26796
rect 7980 26402 8036 30268
rect 8316 30324 8372 30830
rect 8540 30884 8596 30894
rect 8540 30790 8596 30828
rect 8316 30258 8372 30268
rect 8764 30324 8820 30334
rect 8764 30098 8820 30268
rect 8764 30046 8766 30098
rect 8818 30046 8820 30098
rect 8764 30034 8820 30046
rect 8876 29988 8932 30940
rect 9100 30994 9156 31052
rect 9100 30942 9102 30994
rect 9154 30942 9156 30994
rect 9100 30930 9156 30942
rect 9212 30324 9268 31948
rect 9436 31938 9492 31948
rect 9324 31778 9380 31790
rect 9324 31726 9326 31778
rect 9378 31726 9380 31778
rect 9324 31668 9380 31726
rect 9548 31780 9604 32956
rect 9884 32004 9940 32014
rect 9884 31890 9940 31948
rect 9884 31838 9886 31890
rect 9938 31838 9940 31890
rect 9884 31826 9940 31838
rect 10108 31892 10164 31902
rect 10108 31798 10164 31836
rect 9548 31714 9604 31724
rect 9324 31602 9380 31612
rect 9660 31668 9716 31678
rect 9660 31574 9716 31612
rect 9772 31556 9828 31566
rect 9772 31462 9828 31500
rect 10220 31332 10276 34300
rect 10780 33796 10836 38612
rect 11116 38164 11172 38174
rect 11116 38070 11172 38108
rect 10892 37268 10948 37278
rect 10892 37174 10948 37212
rect 11116 36596 11172 36606
rect 11116 36502 11172 36540
rect 11228 36372 11284 45612
rect 11340 45602 11396 45612
rect 12572 45666 12628 45678
rect 12572 45614 12574 45666
rect 12626 45614 12628 45666
rect 11676 45556 11732 45566
rect 11676 45330 11732 45500
rect 11676 45278 11678 45330
rect 11730 45278 11732 45330
rect 11676 45266 11732 45278
rect 12012 45106 12068 45118
rect 12012 45054 12014 45106
rect 12066 45054 12068 45106
rect 11340 44324 11396 44334
rect 11340 44210 11396 44268
rect 11340 44158 11342 44210
rect 11394 44158 11396 44210
rect 11340 44146 11396 44158
rect 11676 44098 11732 44110
rect 11676 44046 11678 44098
rect 11730 44046 11732 44098
rect 11676 43708 11732 44046
rect 11564 43652 11732 43708
rect 12012 43652 12068 45054
rect 12572 43708 12628 45614
rect 12796 45330 12852 45836
rect 13692 45890 13748 45948
rect 14812 46002 15092 46004
rect 14812 45950 14814 46002
rect 14866 45950 15092 46002
rect 14812 45948 15092 45950
rect 16156 46002 16436 46004
rect 16156 45950 16382 46002
rect 16434 45950 16436 46002
rect 16156 45948 16436 45950
rect 14812 45938 14868 45948
rect 13692 45838 13694 45890
rect 13746 45838 13748 45890
rect 13692 45826 13748 45838
rect 15036 45890 15092 45948
rect 15036 45838 15038 45890
rect 15090 45838 15092 45890
rect 15036 45826 15092 45838
rect 16380 45892 16436 45948
rect 16380 45826 16436 45836
rect 17052 45892 17108 45902
rect 17500 45892 17556 49200
rect 18844 46004 18900 49200
rect 20188 46450 20244 49200
rect 20188 46398 20190 46450
rect 20242 46398 20244 46450
rect 18844 46002 19348 46004
rect 18844 45950 18846 46002
rect 18898 45950 19348 46002
rect 18844 45948 19348 45950
rect 18844 45938 18900 45948
rect 17724 45892 17780 45902
rect 17500 45890 17780 45892
rect 17500 45838 17726 45890
rect 17778 45838 17780 45890
rect 17500 45836 17780 45838
rect 17052 45798 17108 45836
rect 12796 45278 12798 45330
rect 12850 45278 12852 45330
rect 12796 45266 12852 45278
rect 14028 45666 14084 45678
rect 14028 45614 14030 45666
rect 14082 45614 14084 45666
rect 12572 43652 12964 43708
rect 11340 43538 11396 43550
rect 11340 43486 11342 43538
rect 11394 43486 11396 43538
rect 11340 43428 11396 43486
rect 11340 43362 11396 43372
rect 11564 42868 11620 43652
rect 12012 43586 12068 43596
rect 12124 43428 12180 43438
rect 11452 42084 11508 42094
rect 11564 42084 11620 42812
rect 11788 43426 12180 43428
rect 11788 43374 12126 43426
rect 12178 43374 12180 43426
rect 11788 43372 12180 43374
rect 11788 42194 11844 43372
rect 12124 43362 12180 43372
rect 12684 42868 12740 42878
rect 12684 42774 12740 42812
rect 11788 42142 11790 42194
rect 11842 42142 11844 42194
rect 11788 42130 11844 42142
rect 11508 42028 11620 42084
rect 11340 41970 11396 41982
rect 11340 41918 11342 41970
rect 11394 41918 11396 41970
rect 11340 41748 11396 41918
rect 11340 41682 11396 41692
rect 11452 38722 11508 42028
rect 11676 41970 11732 41982
rect 11676 41918 11678 41970
rect 11730 41918 11732 41970
rect 11676 41524 11732 41918
rect 11900 41972 11956 41982
rect 11900 41878 11956 41916
rect 11676 41458 11732 41468
rect 12460 41524 12516 41534
rect 11900 41412 11956 41422
rect 11900 41318 11956 41356
rect 12460 41410 12516 41468
rect 12460 41358 12462 41410
rect 12514 41358 12516 41410
rect 12460 41346 12516 41358
rect 12012 41188 12068 41198
rect 12012 41094 12068 41132
rect 12572 41188 12628 41198
rect 12572 41094 12628 41132
rect 11564 41076 11620 41086
rect 11900 41076 11956 41086
rect 11564 41074 11900 41076
rect 11564 41022 11566 41074
rect 11618 41022 11900 41074
rect 11564 41020 11900 41022
rect 11564 41010 11620 41020
rect 11900 40982 11956 41020
rect 12460 40962 12516 40974
rect 12460 40910 12462 40962
rect 12514 40910 12516 40962
rect 12460 40628 12516 40910
rect 12460 40562 12516 40572
rect 12908 40292 12964 43652
rect 13580 42644 13636 42654
rect 13580 42550 13636 42588
rect 13580 41860 13636 41870
rect 13020 41188 13076 41198
rect 13020 40626 13076 41132
rect 13020 40574 13022 40626
rect 13074 40574 13076 40626
rect 13020 40562 13076 40574
rect 13580 40626 13636 41804
rect 13580 40574 13582 40626
rect 13634 40574 13636 40626
rect 13580 40562 13636 40574
rect 13692 40962 13748 40974
rect 13692 40910 13694 40962
rect 13746 40910 13748 40962
rect 13692 40628 13748 40910
rect 13692 40562 13748 40572
rect 13804 40852 13860 40862
rect 13804 40626 13860 40796
rect 13804 40574 13806 40626
rect 13858 40574 13860 40626
rect 13804 40562 13860 40574
rect 13356 40404 13412 40414
rect 13356 40310 13412 40348
rect 13916 40404 13972 40414
rect 13916 40310 13972 40348
rect 12908 40236 13076 40292
rect 12012 39058 12068 39070
rect 12012 39006 12014 39058
rect 12066 39006 12068 39058
rect 11452 38670 11454 38722
rect 11506 38670 11508 38722
rect 11452 38658 11508 38670
rect 11676 38836 11732 38846
rect 11452 37378 11508 37390
rect 11452 37326 11454 37378
rect 11506 37326 11508 37378
rect 11452 36932 11508 37326
rect 11228 36316 11396 36372
rect 10220 31266 10276 31276
rect 10332 33740 10836 33796
rect 10892 36260 10948 36270
rect 10332 31778 10388 33740
rect 10444 33124 10500 33134
rect 10444 32116 10500 33068
rect 10668 32674 10724 32686
rect 10668 32622 10670 32674
rect 10722 32622 10724 32674
rect 10444 32050 10500 32060
rect 10556 32340 10612 32350
rect 10332 31726 10334 31778
rect 10386 31726 10388 31778
rect 9436 31220 9492 31230
rect 9436 31126 9492 31164
rect 9884 31220 9940 31230
rect 9548 30996 9604 31006
rect 9100 30212 9156 30222
rect 9212 30212 9268 30268
rect 9100 30210 9268 30212
rect 9100 30158 9102 30210
rect 9154 30158 9268 30210
rect 9100 30156 9268 30158
rect 9436 30994 9604 30996
rect 9436 30942 9550 30994
rect 9602 30942 9604 30994
rect 9436 30940 9604 30942
rect 9100 30146 9156 30156
rect 9436 30100 9492 30940
rect 9548 30930 9604 30940
rect 9772 30996 9828 31006
rect 9772 30902 9828 30940
rect 9772 30324 9828 30334
rect 9772 30210 9828 30268
rect 9772 30158 9774 30210
rect 9826 30158 9828 30210
rect 9772 30146 9828 30158
rect 8876 29922 8932 29932
rect 9212 30098 9492 30100
rect 9212 30046 9438 30098
rect 9490 30046 9492 30098
rect 9212 30044 9492 30046
rect 9212 29092 9268 30044
rect 9436 30034 9492 30044
rect 8876 29036 9268 29092
rect 8876 28642 8932 29036
rect 8988 28868 9044 28878
rect 8988 28754 9044 28812
rect 8988 28702 8990 28754
rect 9042 28702 9044 28754
rect 8988 28690 9044 28702
rect 8876 28590 8878 28642
rect 8930 28590 8932 28642
rect 8876 28578 8932 28590
rect 9100 28644 9156 28654
rect 9100 28550 9156 28588
rect 8988 28532 9044 28542
rect 8092 27972 8148 27982
rect 8092 27878 8148 27916
rect 8988 27970 9044 28476
rect 9212 28308 9268 29036
rect 9548 28868 9604 28878
rect 9324 28644 9380 28654
rect 9324 28550 9380 28588
rect 9548 28642 9604 28812
rect 9548 28590 9550 28642
rect 9602 28590 9604 28642
rect 9548 28578 9604 28590
rect 9884 28642 9940 31164
rect 9996 30996 10052 31006
rect 10052 30940 10164 30996
rect 9996 30902 10052 30940
rect 10108 30100 10164 30940
rect 10220 30994 10276 31006
rect 10220 30942 10222 30994
rect 10274 30942 10276 30994
rect 10220 30324 10276 30942
rect 10332 30772 10388 31726
rect 10556 30994 10612 32284
rect 10668 32004 10724 32622
rect 10668 31938 10724 31948
rect 10780 31892 10836 31902
rect 10892 31892 10948 36204
rect 11228 36148 11284 36158
rect 11116 36092 11228 36148
rect 11004 32564 11060 32574
rect 11004 32470 11060 32508
rect 10836 31836 10948 31892
rect 10780 31798 10836 31836
rect 11116 31332 11172 36092
rect 11228 36082 11284 36092
rect 10556 30942 10558 30994
rect 10610 30942 10612 30994
rect 10556 30930 10612 30942
rect 10892 31276 11172 31332
rect 11228 31444 11284 31454
rect 10892 31218 10948 31276
rect 10892 31166 10894 31218
rect 10946 31166 10948 31218
rect 10892 30996 10948 31166
rect 10892 30930 10948 30940
rect 10668 30772 10724 30782
rect 10332 30770 10724 30772
rect 10332 30718 10670 30770
rect 10722 30718 10724 30770
rect 10332 30716 10724 30718
rect 10668 30706 10724 30716
rect 10220 30258 10276 30268
rect 10332 30212 10388 30222
rect 10220 30100 10276 30110
rect 10108 30098 10276 30100
rect 10108 30046 10222 30098
rect 10274 30046 10276 30098
rect 10108 30044 10276 30046
rect 10220 29540 10276 30044
rect 9884 28590 9886 28642
rect 9938 28590 9940 28642
rect 9884 28578 9940 28590
rect 9996 28644 10052 28654
rect 9996 28420 10052 28588
rect 10108 28420 10164 28430
rect 9996 28418 10164 28420
rect 9996 28366 10110 28418
rect 10162 28366 10164 28418
rect 9996 28364 10164 28366
rect 9212 28252 9604 28308
rect 9436 28084 9492 28094
rect 9436 27990 9492 28028
rect 8988 27918 8990 27970
rect 9042 27918 9044 27970
rect 8988 27906 9044 27918
rect 9548 27972 9604 28252
rect 9548 27878 9604 27916
rect 8764 27858 8820 27870
rect 8764 27806 8766 27858
rect 8818 27806 8820 27858
rect 8204 27746 8260 27758
rect 8204 27694 8206 27746
rect 8258 27694 8260 27746
rect 8204 27636 8260 27694
rect 8204 27570 8260 27580
rect 8316 27746 8372 27758
rect 8316 27694 8318 27746
rect 8370 27694 8372 27746
rect 8316 27300 8372 27694
rect 8540 27636 8596 27646
rect 8316 27234 8372 27244
rect 8428 27580 8540 27636
rect 7980 26350 7982 26402
rect 8034 26350 8036 26402
rect 7420 25844 7476 25854
rect 7196 25788 7420 25844
rect 6860 25732 6916 25742
rect 6860 25638 6916 25676
rect 6748 25394 6804 25406
rect 6748 25342 6750 25394
rect 6802 25342 6804 25394
rect 6748 23940 6804 25342
rect 6748 23874 6804 23884
rect 7196 23938 7252 25788
rect 7420 25778 7476 25788
rect 7980 25844 8036 26350
rect 8428 26290 8484 27580
rect 8540 27542 8596 27580
rect 8764 26740 8820 27806
rect 8764 26674 8820 26684
rect 8876 27860 8932 27870
rect 8876 26402 8932 27804
rect 9436 27860 9492 27870
rect 8876 26350 8878 26402
rect 8930 26350 8932 26402
rect 8876 26338 8932 26350
rect 9100 26852 9156 26862
rect 8428 26238 8430 26290
rect 8482 26238 8484 26290
rect 8428 26226 8484 26238
rect 8652 26290 8708 26302
rect 8652 26238 8654 26290
rect 8706 26238 8708 26290
rect 8092 26180 8148 26190
rect 8092 26086 8148 26124
rect 8204 26178 8260 26190
rect 8204 26126 8206 26178
rect 8258 26126 8260 26178
rect 7980 25778 8036 25788
rect 8204 25732 8260 26126
rect 8204 25666 8260 25676
rect 8428 26068 8484 26078
rect 7756 25172 7812 25182
rect 7644 24052 7700 24062
rect 7532 23996 7644 24052
rect 7196 23886 7198 23938
rect 7250 23886 7252 23938
rect 6524 23492 6804 23548
rect 6300 22978 6356 22988
rect 5964 22542 5966 22594
rect 6018 22542 6020 22594
rect 5964 22530 6020 22542
rect 4956 22370 5236 22372
rect 4956 22318 4958 22370
rect 5010 22318 5236 22370
rect 4956 22316 5236 22318
rect 4956 22306 5012 22316
rect 4396 21586 4564 21588
rect 4396 21534 4398 21586
rect 4450 21534 4564 21586
rect 4396 21532 4564 21534
rect 5068 21588 5124 22316
rect 5852 22258 5908 22270
rect 5852 22206 5854 22258
rect 5906 22206 5908 22258
rect 5180 21588 5236 21598
rect 5068 21586 5236 21588
rect 5068 21534 5182 21586
rect 5234 21534 5236 21586
rect 5068 21532 5236 21534
rect 4396 21522 4452 21532
rect 5180 21476 5236 21532
rect 5628 21476 5684 21486
rect 5180 21474 5796 21476
rect 5180 21422 5630 21474
rect 5682 21422 5796 21474
rect 5180 21420 5796 21422
rect 5628 21410 5684 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4284 20804 4340 20814
rect 4284 20710 4340 20748
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5068 17780 5124 17790
rect 5068 17686 5124 17724
rect 3948 17154 4004 17164
rect 5740 17442 5796 21420
rect 5852 20804 5908 22206
rect 5852 20738 5908 20748
rect 6636 22260 6692 22270
rect 6524 18452 6580 18462
rect 6524 18358 6580 18396
rect 6636 18338 6692 22204
rect 6636 18286 6638 18338
rect 6690 18286 6692 18338
rect 6076 18228 6132 18238
rect 5740 17390 5742 17442
rect 5794 17390 5796 17442
rect 4060 16996 4116 17006
rect 4060 16902 4116 16940
rect 5740 16884 5796 17390
rect 3164 15428 3220 15438
rect 3164 15334 3220 15372
rect 3500 13748 3556 16492
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5740 16212 5796 16828
rect 5964 18226 6132 18228
rect 5964 18174 6078 18226
rect 6130 18174 6132 18226
rect 5964 18172 6132 18174
rect 5796 16156 5908 16212
rect 5740 16118 5796 16156
rect 5180 15874 5236 15886
rect 5180 15822 5182 15874
rect 5234 15822 5236 15874
rect 5180 15204 5236 15822
rect 5292 15204 5348 15214
rect 5180 15148 5292 15204
rect 5628 15202 5684 15214
rect 5628 15150 5630 15202
rect 5682 15150 5684 15202
rect 5628 15148 5684 15150
rect 5292 15110 5348 15148
rect 5404 15092 5684 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 3500 13682 3556 13692
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 5404 11844 5460 15092
rect 5852 14642 5908 16156
rect 5964 15988 6020 18172
rect 6076 18162 6132 18172
rect 6636 17892 6692 18286
rect 6188 17836 6692 17892
rect 6188 17780 6244 17836
rect 6748 17780 6804 23492
rect 7084 23268 7140 23278
rect 7196 23268 7252 23886
rect 7420 23938 7476 23950
rect 7420 23886 7422 23938
rect 7474 23886 7476 23938
rect 7420 23604 7476 23886
rect 7420 23538 7476 23548
rect 7084 23266 7252 23268
rect 7084 23214 7086 23266
rect 7138 23214 7252 23266
rect 7084 23212 7252 23214
rect 7084 23202 7140 23212
rect 7308 23156 7364 23166
rect 7308 23062 7364 23100
rect 7532 23154 7588 23996
rect 7644 23958 7700 23996
rect 7532 23102 7534 23154
rect 7586 23102 7588 23154
rect 7196 23042 7252 23054
rect 7196 22990 7198 23042
rect 7250 22990 7252 23042
rect 6076 17554 6132 17566
rect 6076 17502 6078 17554
rect 6130 17502 6132 17554
rect 6076 16884 6132 17502
rect 6188 17554 6244 17724
rect 6188 17502 6190 17554
rect 6242 17502 6244 17554
rect 6188 17490 6244 17502
rect 6300 17724 6804 17780
rect 7084 22820 7140 22830
rect 6076 16098 6132 16828
rect 6188 16772 6244 16782
rect 6188 16678 6244 16716
rect 6076 16046 6078 16098
rect 6130 16046 6132 16098
rect 6076 16034 6132 16046
rect 5964 15922 6020 15932
rect 6188 15988 6244 15998
rect 6300 15988 6356 17724
rect 6412 17556 6468 17566
rect 6636 17556 6692 17566
rect 6412 17554 6692 17556
rect 6412 17502 6414 17554
rect 6466 17502 6638 17554
rect 6690 17502 6692 17554
rect 6412 17500 6692 17502
rect 6412 17490 6468 17500
rect 6636 17490 6692 17500
rect 6748 17556 6804 17566
rect 6748 17462 6804 17500
rect 6972 17556 7028 17566
rect 6972 17462 7028 17500
rect 7084 17332 7140 22764
rect 7196 22484 7252 22990
rect 7196 22418 7252 22428
rect 7532 22148 7588 23102
rect 7644 23714 7700 23726
rect 7644 23662 7646 23714
rect 7698 23662 7700 23714
rect 7644 22596 7700 23662
rect 7756 23492 7812 25116
rect 8204 24836 8260 24846
rect 7868 23940 7924 23950
rect 7868 23846 7924 23884
rect 8204 23938 8260 24780
rect 8204 23886 8206 23938
rect 8258 23886 8260 23938
rect 8204 23874 8260 23886
rect 7756 23436 7924 23492
rect 7756 23154 7812 23166
rect 7756 23102 7758 23154
rect 7810 23102 7812 23154
rect 7756 23044 7812 23102
rect 7756 22978 7812 22988
rect 7644 22530 7700 22540
rect 7532 22082 7588 22092
rect 7644 21476 7700 21486
rect 7644 21382 7700 21420
rect 7196 19124 7252 19134
rect 7196 18452 7252 19068
rect 7196 18358 7252 18396
rect 7644 18338 7700 18350
rect 7644 18286 7646 18338
rect 7698 18286 7700 18338
rect 6972 17276 7140 17332
rect 7196 18226 7252 18238
rect 7196 18174 7198 18226
rect 7250 18174 7252 18226
rect 7196 17666 7252 18174
rect 7644 18226 7700 18286
rect 7644 18174 7646 18226
rect 7698 18174 7700 18226
rect 7644 18162 7700 18174
rect 7868 18340 7924 23436
rect 7980 23156 8036 23166
rect 7980 23062 8036 23100
rect 8316 23044 8372 23054
rect 8316 22950 8372 22988
rect 8316 22148 8372 22158
rect 8316 22054 8372 22092
rect 8428 21812 8484 26012
rect 8652 25284 8708 26238
rect 8652 25218 8708 25228
rect 8988 24836 9044 24846
rect 8876 24500 8932 24510
rect 8764 24052 8820 24062
rect 8652 23996 8764 24052
rect 8540 23716 8596 23726
rect 8652 23716 8708 23996
rect 8764 23986 8820 23996
rect 8540 23714 8708 23716
rect 8540 23662 8542 23714
rect 8594 23662 8708 23714
rect 8540 23660 8708 23662
rect 8540 23650 8596 23660
rect 8876 23154 8932 24444
rect 8876 23102 8878 23154
rect 8930 23102 8932 23154
rect 8876 23090 8932 23102
rect 8652 23044 8708 23054
rect 8652 23042 8820 23044
rect 8652 22990 8654 23042
rect 8706 22990 8820 23042
rect 8652 22988 8820 22990
rect 8652 22978 8708 22988
rect 8764 22484 8820 22988
rect 8764 22428 8932 22484
rect 8764 22260 8820 22270
rect 8764 22166 8820 22204
rect 8876 22148 8932 22428
rect 8988 22370 9044 24780
rect 9100 22708 9156 26796
rect 9436 22820 9492 27804
rect 9772 27748 9828 27758
rect 9772 27654 9828 27692
rect 9996 27746 10052 28364
rect 10108 28354 10164 28364
rect 10220 28084 10276 29484
rect 9996 27694 9998 27746
rect 10050 27694 10052 27746
rect 9884 27636 9940 27646
rect 9996 27636 10052 27694
rect 9940 27580 10052 27636
rect 10108 28028 10276 28084
rect 9884 27570 9940 27580
rect 10108 27524 10164 28028
rect 10332 27972 10388 30156
rect 10444 28532 10500 28542
rect 11228 28532 11284 31388
rect 11340 30100 11396 36316
rect 11452 36036 11508 36876
rect 11564 36820 11620 36830
rect 11564 36482 11620 36764
rect 11564 36430 11566 36482
rect 11618 36430 11620 36482
rect 11564 36418 11620 36430
rect 11676 36148 11732 38780
rect 11900 38724 11956 38734
rect 11788 38668 11900 38724
rect 11788 37044 11844 38668
rect 11900 38630 11956 38668
rect 11900 38500 11956 38510
rect 11900 37490 11956 38444
rect 11900 37438 11902 37490
rect 11954 37438 11956 37490
rect 11900 37426 11956 37438
rect 12012 37268 12068 39006
rect 12572 39060 12628 39070
rect 12572 38966 12628 39004
rect 12460 38948 12516 38958
rect 12124 38836 12180 38846
rect 12124 38742 12180 38780
rect 12460 38834 12516 38892
rect 12460 38782 12462 38834
rect 12514 38782 12516 38834
rect 12460 38770 12516 38782
rect 12796 38834 12852 38846
rect 12796 38782 12798 38834
rect 12850 38782 12852 38834
rect 12460 38500 12516 38510
rect 12460 38162 12516 38444
rect 12460 38110 12462 38162
rect 12514 38110 12516 38162
rect 12460 38098 12516 38110
rect 12460 37380 12516 37390
rect 12460 37286 12516 37324
rect 12796 37380 12852 38782
rect 12796 37314 12852 37324
rect 12012 37202 12068 37212
rect 12572 37268 12628 37278
rect 12460 37044 12516 37054
rect 11788 36988 12292 37044
rect 12012 36708 12068 36718
rect 12012 36614 12068 36652
rect 12236 36596 12292 36988
rect 12236 36502 12292 36540
rect 12460 36482 12516 36988
rect 12460 36430 12462 36482
rect 12514 36430 12516 36482
rect 12460 36418 12516 36430
rect 11788 36372 11844 36382
rect 11788 36278 11844 36316
rect 12012 36260 12068 36270
rect 12012 36258 12180 36260
rect 12012 36206 12014 36258
rect 12066 36206 12180 36258
rect 12012 36204 12180 36206
rect 12012 36194 12068 36204
rect 11676 36082 11732 36092
rect 11564 36036 11620 36046
rect 11452 35980 11564 36036
rect 11564 35970 11620 35980
rect 11676 35924 11732 35934
rect 11676 35028 11732 35868
rect 12012 35474 12068 35486
rect 12012 35422 12014 35474
rect 12066 35422 12068 35474
rect 12012 35140 12068 35422
rect 11900 35084 12068 35140
rect 12124 35140 12180 36204
rect 11676 34972 11788 35028
rect 11732 34916 11788 34972
rect 11732 34860 11844 34916
rect 11788 34580 11844 34860
rect 11788 34514 11844 34524
rect 11564 33906 11620 33918
rect 11564 33854 11566 33906
rect 11618 33854 11620 33906
rect 11452 31554 11508 31566
rect 11452 31502 11454 31554
rect 11506 31502 11508 31554
rect 11452 31108 11508 31502
rect 11564 31220 11620 33854
rect 11900 31892 11956 35084
rect 12124 35074 12180 35084
rect 12236 36148 12292 36158
rect 12460 36148 12516 36158
rect 12236 34914 12292 36092
rect 12348 36092 12460 36148
rect 12348 35698 12404 36092
rect 12460 36082 12516 36092
rect 12348 35646 12350 35698
rect 12402 35646 12404 35698
rect 12348 35634 12404 35646
rect 12572 35586 12628 37212
rect 12684 37266 12740 37278
rect 12684 37214 12686 37266
rect 12738 37214 12740 37266
rect 12684 37156 12740 37214
rect 12684 37090 12740 37100
rect 12908 36484 12964 36494
rect 12572 35534 12574 35586
rect 12626 35534 12628 35586
rect 12572 35522 12628 35534
rect 12684 36372 12740 36382
rect 12236 34862 12238 34914
rect 12290 34862 12292 34914
rect 12236 34850 12292 34862
rect 12348 35364 12404 35374
rect 12684 35308 12740 36316
rect 12236 34580 12292 34590
rect 12236 34242 12292 34524
rect 12236 34190 12238 34242
rect 12290 34190 12292 34242
rect 12236 34178 12292 34190
rect 12348 34242 12404 35308
rect 12572 35252 12740 35308
rect 12908 36258 12964 36428
rect 12908 36206 12910 36258
rect 12962 36206 12964 36258
rect 12572 35028 12628 35252
rect 12460 34972 12628 35028
rect 12460 34690 12516 34972
rect 12572 34804 12628 34814
rect 12572 34710 12628 34748
rect 12908 34804 12964 36206
rect 12908 34738 12964 34748
rect 12460 34638 12462 34690
rect 12514 34638 12516 34690
rect 12460 34356 12516 34638
rect 12684 34690 12740 34702
rect 12684 34638 12686 34690
rect 12738 34638 12740 34690
rect 12684 34356 12740 34638
rect 12460 34300 12628 34356
rect 12348 34190 12350 34242
rect 12402 34190 12404 34242
rect 12348 34178 12404 34190
rect 12012 34130 12068 34142
rect 12012 34078 12014 34130
rect 12066 34078 12068 34130
rect 12012 33460 12068 34078
rect 12012 33394 12068 33404
rect 12460 34130 12516 34142
rect 12460 34078 12462 34130
rect 12514 34078 12516 34130
rect 12460 33124 12516 34078
rect 12012 33068 12516 33124
rect 12012 32786 12068 33068
rect 12012 32734 12014 32786
rect 12066 32734 12068 32786
rect 12012 32722 12068 32734
rect 11564 31154 11620 31164
rect 11788 31836 11956 31892
rect 12348 32676 12404 32686
rect 12572 32676 12628 34300
rect 12684 34290 12740 34300
rect 12796 34690 12852 34702
rect 12796 34638 12798 34690
rect 12850 34638 12852 34690
rect 12796 33348 12852 34638
rect 12796 33282 12852 33292
rect 12908 33124 12964 33134
rect 12796 33122 12964 33124
rect 12796 33070 12910 33122
rect 12962 33070 12964 33122
rect 12796 33068 12964 33070
rect 12684 32676 12740 32686
rect 12572 32620 12684 32676
rect 12348 32562 12404 32620
rect 12684 32610 12740 32620
rect 12348 32510 12350 32562
rect 12402 32510 12404 32562
rect 11452 31042 11508 31052
rect 11452 30882 11508 30894
rect 11452 30830 11454 30882
rect 11506 30830 11508 30882
rect 11452 30770 11508 30830
rect 11452 30718 11454 30770
rect 11506 30718 11508 30770
rect 11452 30706 11508 30718
rect 11788 30212 11844 31836
rect 12124 31780 12180 31790
rect 12124 31686 12180 31724
rect 11900 31666 11956 31678
rect 11900 31614 11902 31666
rect 11954 31614 11956 31666
rect 11900 30996 11956 31614
rect 11900 30930 11956 30940
rect 12012 31666 12068 31678
rect 12012 31614 12014 31666
rect 12066 31614 12068 31666
rect 11788 30146 11844 30156
rect 11340 30034 11396 30044
rect 11788 29540 11844 29550
rect 11676 29484 11788 29540
rect 11340 28532 11396 28542
rect 10444 28530 10836 28532
rect 10444 28478 10446 28530
rect 10498 28478 10836 28530
rect 10444 28476 10836 28478
rect 11228 28476 11340 28532
rect 10444 28466 10500 28476
rect 10780 28082 10836 28476
rect 10780 28030 10782 28082
rect 10834 28030 10836 28082
rect 10444 27972 10500 27982
rect 10332 27970 10500 27972
rect 10332 27918 10446 27970
rect 10498 27918 10500 27970
rect 10332 27916 10500 27918
rect 10444 27906 10500 27916
rect 9996 27468 10164 27524
rect 10220 27858 10276 27870
rect 10220 27806 10222 27858
rect 10274 27806 10276 27858
rect 9996 27412 10052 27468
rect 9884 27356 10052 27412
rect 9884 27186 9940 27356
rect 9884 27134 9886 27186
rect 9938 27134 9940 27186
rect 9884 27122 9940 27134
rect 9996 27076 10052 27086
rect 9772 26402 9828 26414
rect 9772 26350 9774 26402
rect 9826 26350 9828 26402
rect 9772 24052 9828 26350
rect 9996 26290 10052 27020
rect 10220 26852 10276 27806
rect 10444 27076 10500 27086
rect 10780 27076 10836 28030
rect 11340 27858 11396 28476
rect 11340 27806 11342 27858
rect 11394 27806 11396 27858
rect 11340 27794 11396 27806
rect 11564 27412 11620 27422
rect 11564 27188 11620 27356
rect 10500 27020 10836 27076
rect 10444 26982 10500 27020
rect 10780 26962 10836 27020
rect 10780 26910 10782 26962
rect 10834 26910 10836 26962
rect 10780 26898 10836 26910
rect 11116 27186 11620 27188
rect 11116 27134 11566 27186
rect 11618 27134 11620 27186
rect 11116 27132 11620 27134
rect 11116 27074 11172 27132
rect 11564 27122 11620 27132
rect 11116 27022 11118 27074
rect 11170 27022 11172 27074
rect 11116 26908 11172 27022
rect 10220 26786 10276 26796
rect 11004 26852 11172 26908
rect 9996 26238 9998 26290
rect 10050 26238 10052 26290
rect 9996 26226 10052 26238
rect 9996 26068 10052 26078
rect 9772 23986 9828 23996
rect 9884 24612 9940 24622
rect 9436 22754 9492 22764
rect 9772 23042 9828 23054
rect 9772 22990 9774 23042
rect 9826 22990 9828 23042
rect 9100 22642 9156 22652
rect 9772 22484 9828 22990
rect 8988 22318 8990 22370
rect 9042 22318 9044 22370
rect 8988 22306 9044 22318
rect 9212 22428 9828 22484
rect 9884 22482 9940 24556
rect 9884 22430 9886 22482
rect 9938 22430 9940 22482
rect 9100 22148 9156 22158
rect 8876 22146 9156 22148
rect 8876 22094 9102 22146
rect 9154 22094 9156 22146
rect 8876 22092 9156 22094
rect 9100 22082 9156 22092
rect 9212 22146 9268 22428
rect 9884 22260 9940 22430
rect 9996 22484 10052 26012
rect 10668 26068 10724 26078
rect 10668 23940 10724 26012
rect 10668 23874 10724 23884
rect 9996 22428 10164 22484
rect 9660 22204 9940 22260
rect 9996 22260 10052 22270
rect 9212 22094 9214 22146
rect 9266 22094 9268 22146
rect 8428 21756 8596 21812
rect 8428 21586 8484 21598
rect 8428 21534 8430 21586
rect 8482 21534 8484 21586
rect 8092 21474 8148 21486
rect 8092 21422 8094 21474
rect 8146 21422 8148 21474
rect 8092 20580 8148 21422
rect 8428 21476 8484 21534
rect 8316 20580 8372 20590
rect 8092 20524 8316 20580
rect 7980 19908 8036 19918
rect 7980 19814 8036 19852
rect 8316 19906 8372 20524
rect 8316 19854 8318 19906
rect 8370 19854 8372 19906
rect 8316 19236 8372 19854
rect 8428 19684 8484 21420
rect 8428 19618 8484 19628
rect 8316 19170 8372 19180
rect 8540 18788 8596 21756
rect 8988 21700 9044 21710
rect 8988 21606 9044 21644
rect 8988 21252 9044 21262
rect 8988 20130 9044 21196
rect 9100 20580 9156 20590
rect 9100 20486 9156 20524
rect 8988 20078 8990 20130
rect 9042 20078 9044 20130
rect 8988 20066 9044 20078
rect 9212 20132 9268 22094
rect 9324 22148 9380 22158
rect 9660 22148 9716 22204
rect 9324 22146 9716 22148
rect 9324 22094 9326 22146
rect 9378 22094 9716 22146
rect 9324 22092 9716 22094
rect 9324 22082 9380 22092
rect 9548 21588 9604 21598
rect 9436 21586 9604 21588
rect 9436 21534 9550 21586
rect 9602 21534 9604 21586
rect 9436 21532 9604 21534
rect 9436 20580 9492 21532
rect 9548 21522 9604 21532
rect 9660 21588 9716 21598
rect 9660 21494 9716 21532
rect 9996 20914 10052 22204
rect 10108 22036 10164 22428
rect 10108 21970 10164 21980
rect 10668 22370 10724 22382
rect 10668 22318 10670 22370
rect 10722 22318 10724 22370
rect 10108 21698 10164 21710
rect 10108 21646 10110 21698
rect 10162 21646 10164 21698
rect 10108 21588 10164 21646
rect 10668 21588 10724 22318
rect 10164 21532 10388 21588
rect 10108 21522 10164 21532
rect 9996 20862 9998 20914
rect 10050 20862 10052 20914
rect 9996 20850 10052 20862
rect 10332 20802 10388 21532
rect 10668 21522 10724 21532
rect 11004 21028 11060 26852
rect 11676 24834 11732 29484
rect 11788 29474 11844 29484
rect 12012 25620 12068 31614
rect 12348 29540 12404 32510
rect 12460 32564 12516 32574
rect 12460 32004 12516 32508
rect 12572 32452 12628 32462
rect 12796 32452 12852 33068
rect 12908 33058 12964 33068
rect 12908 32564 12964 32574
rect 12908 32470 12964 32508
rect 12572 32450 12852 32452
rect 12572 32398 12574 32450
rect 12626 32398 12852 32450
rect 12572 32396 12852 32398
rect 12572 32386 12628 32396
rect 12572 32004 12628 32014
rect 12460 32002 12628 32004
rect 12460 31950 12574 32002
rect 12626 31950 12628 32002
rect 12460 31948 12628 31950
rect 12572 31938 12628 31948
rect 12684 31666 12740 32396
rect 12684 31614 12686 31666
rect 12738 31614 12740 31666
rect 12684 31556 12740 31614
rect 12684 31490 12740 31500
rect 13020 30212 13076 40236
rect 13916 39956 13972 39966
rect 13692 39620 13748 39630
rect 13468 38948 13524 38958
rect 13468 38724 13524 38892
rect 13692 38836 13748 39564
rect 13916 39060 13972 39900
rect 13916 38966 13972 39004
rect 13580 38724 13636 38734
rect 13468 38722 13636 38724
rect 13468 38670 13582 38722
rect 13634 38670 13636 38722
rect 13468 38668 13636 38670
rect 13244 37156 13300 37166
rect 13244 37062 13300 37100
rect 13356 36708 13412 36718
rect 13132 36596 13188 36606
rect 13132 35364 13188 36540
rect 13132 35298 13188 35308
rect 13356 35588 13412 36652
rect 13468 36484 13524 38668
rect 13580 38658 13636 38668
rect 13692 38162 13748 38780
rect 13692 38110 13694 38162
rect 13746 38110 13748 38162
rect 13692 38098 13748 38110
rect 13916 38052 13972 38062
rect 13804 37492 13860 37502
rect 13804 37398 13860 37436
rect 13916 36708 13972 37996
rect 14028 36932 14084 45614
rect 15260 45668 15316 45678
rect 14700 45220 14756 45230
rect 14700 44322 14756 45164
rect 15260 44434 15316 45612
rect 15260 44382 15262 44434
rect 15314 44382 15316 44434
rect 15260 44370 15316 44382
rect 15372 45666 15428 45678
rect 15372 45614 15374 45666
rect 15426 45614 15428 45666
rect 14700 44270 14702 44322
rect 14754 44270 14756 44322
rect 14700 44258 14756 44270
rect 14812 44100 14868 44110
rect 14812 44006 14868 44044
rect 15148 44100 15204 44110
rect 15148 44006 15204 44044
rect 14252 43652 14308 43662
rect 14252 43426 14308 43596
rect 14252 43374 14254 43426
rect 14306 43374 14308 43426
rect 14252 39620 14308 43374
rect 14812 43428 14868 43438
rect 14812 43334 14868 43372
rect 15036 42866 15092 42878
rect 15036 42814 15038 42866
rect 15090 42814 15092 42866
rect 14700 42084 14756 42094
rect 14364 40852 14420 40862
rect 14364 40626 14420 40796
rect 14364 40574 14366 40626
rect 14418 40574 14420 40626
rect 14364 40562 14420 40574
rect 14252 39564 14532 39620
rect 14140 39396 14196 39406
rect 14140 39302 14196 39340
rect 14252 39394 14308 39406
rect 14252 39342 14254 39394
rect 14306 39342 14308 39394
rect 14252 39284 14308 39342
rect 14252 39218 14308 39228
rect 14364 39172 14420 39182
rect 14364 38388 14420 39116
rect 14476 39058 14532 39564
rect 14476 39006 14478 39058
rect 14530 39006 14532 39058
rect 14476 38994 14532 39006
rect 14588 39618 14644 39630
rect 14588 39566 14590 39618
rect 14642 39566 14644 39618
rect 14588 38836 14644 39566
rect 14700 39506 14756 42028
rect 15036 42084 15092 42814
rect 15036 42018 15092 42028
rect 15036 39732 15092 39742
rect 15036 39638 15092 39676
rect 15372 39730 15428 45614
rect 17276 45666 17332 45678
rect 17276 45614 17278 45666
rect 17330 45614 17332 45666
rect 16380 44434 16436 44446
rect 16380 44382 16382 44434
rect 16434 44382 16436 44434
rect 16380 43652 16436 44382
rect 15372 39678 15374 39730
rect 15426 39678 15428 39730
rect 15372 39666 15428 39678
rect 15484 42532 15540 42542
rect 14700 39454 14702 39506
rect 14754 39454 14756 39506
rect 14700 39172 14756 39454
rect 14700 39106 14756 39116
rect 14812 39394 14868 39406
rect 14812 39342 14814 39394
rect 14866 39342 14868 39394
rect 14588 38770 14644 38780
rect 14700 38946 14756 38958
rect 14700 38894 14702 38946
rect 14754 38894 14756 38946
rect 14700 38724 14756 38894
rect 14364 38322 14420 38332
rect 14476 38612 14756 38668
rect 14476 38052 14532 38612
rect 14252 37996 14532 38052
rect 14252 37378 14308 37996
rect 14812 37492 14868 39342
rect 15036 38836 15092 38846
rect 15036 38724 15092 38780
rect 15260 38834 15316 38846
rect 15260 38782 15262 38834
rect 15314 38782 15316 38834
rect 15260 38724 15316 38782
rect 15036 38668 15316 38724
rect 15484 38668 15540 42476
rect 16380 42532 16436 43596
rect 17276 42868 17332 45614
rect 17612 45330 17668 45836
rect 17724 45826 17780 45836
rect 19292 45890 19348 45948
rect 20188 46002 20244 46398
rect 20188 45950 20190 46002
rect 20242 45950 20244 46002
rect 20188 45938 20244 45950
rect 20972 46450 21028 46462
rect 20972 46398 20974 46450
rect 21026 46398 21028 46450
rect 19292 45838 19294 45890
rect 19346 45838 19348 45890
rect 19292 45826 19348 45838
rect 20972 45890 21028 46398
rect 20972 45838 20974 45890
rect 21026 45838 21028 45890
rect 20972 45826 21028 45838
rect 21532 46116 21588 49200
rect 21532 46060 22036 46116
rect 18956 45780 19012 45790
rect 18060 45668 18116 45678
rect 18060 45666 18228 45668
rect 18060 45614 18062 45666
rect 18114 45614 18228 45666
rect 18060 45612 18228 45614
rect 18060 45602 18116 45612
rect 17612 45278 17614 45330
rect 17666 45278 17668 45330
rect 17612 45266 17668 45278
rect 17948 43652 18004 43662
rect 17948 43558 18004 43596
rect 18060 43538 18116 43550
rect 18060 43486 18062 43538
rect 18114 43486 18116 43538
rect 17052 42812 17276 42868
rect 16380 42466 16436 42476
rect 16604 42644 16660 42654
rect 16380 40404 16436 40414
rect 14252 37326 14254 37378
rect 14306 37326 14308 37378
rect 14252 37314 14308 37326
rect 14364 37436 14868 37492
rect 14924 38612 15092 38668
rect 15372 38612 15540 38668
rect 15708 39732 15764 39742
rect 14028 36866 14084 36876
rect 13692 36652 13972 36708
rect 13580 36596 13636 36634
rect 13580 36530 13636 36540
rect 13468 36260 13524 36428
rect 13692 36482 13748 36652
rect 14028 36596 14084 36606
rect 13692 36430 13694 36482
rect 13746 36430 13748 36482
rect 13692 36372 13748 36430
rect 13468 36194 13524 36204
rect 13580 36316 13748 36372
rect 13916 36482 13972 36494
rect 13916 36430 13918 36482
rect 13970 36430 13972 36482
rect 13580 35700 13636 36316
rect 13916 36260 13972 36430
rect 14028 36482 14084 36540
rect 14028 36430 14030 36482
rect 14082 36430 14084 36482
rect 14028 36418 14084 36430
rect 14364 36372 14420 37436
rect 14812 37268 14868 37278
rect 14924 37268 14980 38612
rect 14812 37266 14980 37268
rect 14812 37214 14814 37266
rect 14866 37214 14980 37266
rect 14812 37212 14980 37214
rect 15372 37266 15428 38612
rect 15372 37214 15374 37266
rect 15426 37214 15428 37266
rect 14812 37202 14868 37212
rect 15372 37202 15428 37214
rect 13916 36194 13972 36204
rect 14252 36316 14420 36372
rect 14476 37154 14532 37166
rect 14476 37102 14478 37154
rect 14530 37102 14532 37154
rect 14028 35700 14084 35710
rect 13580 35698 14084 35700
rect 13580 35646 14030 35698
rect 14082 35646 14084 35698
rect 13580 35644 14084 35646
rect 14028 35634 14084 35644
rect 13132 34356 13188 34366
rect 13132 34262 13188 34300
rect 13244 32788 13300 32798
rect 13356 32788 13412 35532
rect 14028 35140 14084 35150
rect 13692 35028 13748 35038
rect 13692 34934 13748 34972
rect 13468 34916 13524 34926
rect 13468 34354 13524 34860
rect 13468 34302 13470 34354
rect 13522 34302 13524 34354
rect 13468 34290 13524 34302
rect 14028 34242 14084 35084
rect 14028 34190 14030 34242
rect 14082 34190 14084 34242
rect 14028 34178 14084 34190
rect 13244 32786 13412 32788
rect 13244 32734 13246 32786
rect 13298 32734 13412 32786
rect 13244 32732 13412 32734
rect 13244 32722 13300 32732
rect 13356 31780 13412 32732
rect 13916 34130 13972 34142
rect 13916 34078 13918 34130
rect 13970 34078 13972 34130
rect 13356 31714 13412 31724
rect 13692 32676 13748 32686
rect 13692 32564 13748 32620
rect 13804 32564 13860 32574
rect 13692 32562 13860 32564
rect 13692 32510 13806 32562
rect 13858 32510 13860 32562
rect 13692 32508 13860 32510
rect 13468 31556 13524 31566
rect 13580 31556 13636 31566
rect 13524 31554 13636 31556
rect 13524 31502 13582 31554
rect 13634 31502 13636 31554
rect 13524 31500 13636 31502
rect 13244 30882 13300 30894
rect 13244 30830 13246 30882
rect 13298 30830 13300 30882
rect 13244 30436 13300 30830
rect 13468 30548 13524 31500
rect 13580 31490 13636 31500
rect 13468 30482 13524 30492
rect 13580 30994 13636 31006
rect 13580 30942 13582 30994
rect 13634 30942 13636 30994
rect 13244 30370 13300 30380
rect 13580 30436 13636 30942
rect 13580 30370 13636 30380
rect 13692 30212 13748 32508
rect 13804 32498 13860 32508
rect 13916 31892 13972 34078
rect 14252 34130 14308 36316
rect 14364 35700 14420 35710
rect 14364 35606 14420 35644
rect 14476 34580 14532 37102
rect 15148 37156 15204 37166
rect 14812 36932 14868 36942
rect 14868 36876 14980 36932
rect 14812 36866 14868 36876
rect 14812 36484 14868 36494
rect 14700 36258 14756 36270
rect 14700 36206 14702 36258
rect 14754 36206 14756 36258
rect 14700 35924 14756 36206
rect 14700 35858 14756 35868
rect 14812 36260 14868 36428
rect 14812 35922 14868 36204
rect 14812 35870 14814 35922
rect 14866 35870 14868 35922
rect 14812 35858 14868 35870
rect 14476 34514 14532 34524
rect 14252 34078 14254 34130
rect 14306 34078 14308 34130
rect 14252 34066 14308 34078
rect 14364 32564 14420 32574
rect 14364 32470 14420 32508
rect 14924 31892 14980 36876
rect 15148 36482 15204 37100
rect 15596 36596 15652 36606
rect 15596 36502 15652 36540
rect 15148 36430 15150 36482
rect 15202 36430 15204 36482
rect 13916 31826 13972 31836
rect 14476 31890 14980 31892
rect 14476 31838 14926 31890
rect 14978 31838 14980 31890
rect 14476 31836 14980 31838
rect 14028 31780 14084 31790
rect 13020 30146 13076 30156
rect 13580 30156 13748 30212
rect 13804 31668 13860 31678
rect 13804 31106 13860 31612
rect 13804 31054 13806 31106
rect 13858 31054 13860 31106
rect 12348 29474 12404 29484
rect 13132 30100 13188 30110
rect 13132 28420 13188 30044
rect 13580 29316 13636 30156
rect 13692 29540 13748 29550
rect 13692 29446 13748 29484
rect 13580 29260 13748 29316
rect 13692 28868 13748 29260
rect 13804 28980 13860 31054
rect 14028 30994 14084 31724
rect 14028 30942 14030 30994
rect 14082 30942 14084 30994
rect 14028 30930 14084 30942
rect 14476 31106 14532 31836
rect 14924 31826 14980 31836
rect 15036 35924 15092 35934
rect 14588 31220 14644 31230
rect 14588 31126 14644 31164
rect 14476 31054 14478 31106
rect 14530 31054 14532 31106
rect 14252 30884 14308 30894
rect 14252 30790 14308 30828
rect 14476 30884 14532 31054
rect 14476 30818 14532 30828
rect 14812 30772 14868 30782
rect 14812 30678 14868 30716
rect 14028 30548 14084 30558
rect 13916 30324 13972 30334
rect 13916 29092 13972 30268
rect 14028 29426 14084 30492
rect 15036 30436 15092 35868
rect 15036 30370 15092 30380
rect 15148 35588 15204 36430
rect 15484 36484 15540 36494
rect 15484 36260 15540 36428
rect 15484 36194 15540 36204
rect 15708 36484 15764 39676
rect 16044 39732 16100 39742
rect 16044 38834 16100 39676
rect 16044 38782 16046 38834
rect 16098 38782 16100 38834
rect 16044 38770 16100 38782
rect 16156 39396 16212 39406
rect 16156 37378 16212 39340
rect 16268 39394 16324 39406
rect 16268 39342 16270 39394
rect 16322 39342 16324 39394
rect 16268 39172 16324 39342
rect 16268 39106 16324 39116
rect 16380 38668 16436 40348
rect 16492 39060 16548 39070
rect 16492 38834 16548 39004
rect 16492 38782 16494 38834
rect 16546 38782 16548 38834
rect 16492 38770 16548 38782
rect 16156 37326 16158 37378
rect 16210 37326 16212 37378
rect 15820 37268 15876 37278
rect 15820 37174 15876 37212
rect 16156 36596 16212 37326
rect 15708 36428 16100 36484
rect 15708 35924 15764 36428
rect 15708 35830 15764 35868
rect 15932 36258 15988 36270
rect 15932 36206 15934 36258
rect 15986 36206 15988 36258
rect 15260 35588 15316 35598
rect 15148 35586 15316 35588
rect 15148 35534 15262 35586
rect 15314 35534 15316 35586
rect 15148 35532 15316 35534
rect 15148 30324 15204 35532
rect 15260 35522 15316 35532
rect 15932 35252 15988 36206
rect 16044 36260 16100 36428
rect 16156 36370 16212 36540
rect 16156 36318 16158 36370
rect 16210 36318 16212 36370
rect 16156 36306 16212 36318
rect 16268 38612 16436 38668
rect 16044 35922 16100 36204
rect 16044 35870 16046 35922
rect 16098 35870 16100 35922
rect 16044 35858 16100 35870
rect 15932 35186 15988 35196
rect 15372 34580 15428 34590
rect 15260 31108 15316 31118
rect 15260 31014 15316 31052
rect 15372 31106 15428 34524
rect 15596 32564 15652 32574
rect 15372 31054 15374 31106
rect 15426 31054 15428 31106
rect 15372 31042 15428 31054
rect 15484 32508 15596 32564
rect 15148 30268 15316 30324
rect 14252 30212 14308 30222
rect 14252 30118 14308 30156
rect 14700 30212 14756 30222
rect 14700 30118 14756 30156
rect 15036 30212 15092 30222
rect 14476 29988 14532 29998
rect 14476 29894 14532 29932
rect 14028 29374 14030 29426
rect 14082 29374 14084 29426
rect 14028 29316 14084 29374
rect 14812 29876 14868 29886
rect 14812 29426 14868 29820
rect 14812 29374 14814 29426
rect 14866 29374 14868 29426
rect 14812 29362 14868 29374
rect 14028 29260 14308 29316
rect 13916 29036 14196 29092
rect 13804 28924 13972 28980
rect 13692 28812 13860 28868
rect 13132 28354 13188 28364
rect 13692 28308 13748 28318
rect 12012 25554 12068 25564
rect 13020 26516 13076 26526
rect 11676 24782 11678 24834
rect 11730 24782 11732 24834
rect 11116 24724 11172 24734
rect 11116 22482 11172 24668
rect 11676 24500 11732 24782
rect 11788 24724 11844 24734
rect 11788 24630 11844 24668
rect 12236 24724 12292 24734
rect 11676 24434 11732 24444
rect 11900 24610 11956 24622
rect 11900 24558 11902 24610
rect 11954 24558 11956 24610
rect 11564 23996 11844 24052
rect 11564 23938 11620 23996
rect 11564 23886 11566 23938
rect 11618 23886 11620 23938
rect 11564 23874 11620 23886
rect 11676 23828 11732 23838
rect 11676 23380 11732 23772
rect 11116 22430 11118 22482
rect 11170 22430 11172 22482
rect 11116 22418 11172 22430
rect 11564 23324 11732 23380
rect 11452 21812 11508 21822
rect 11452 21718 11508 21756
rect 11564 21700 11620 23324
rect 11676 23154 11732 23166
rect 11676 23102 11678 23154
rect 11730 23102 11732 23154
rect 11676 22372 11732 23102
rect 11788 22484 11844 23996
rect 11900 23828 11956 24558
rect 12236 23940 12292 24668
rect 12460 24722 12516 24734
rect 12460 24670 12462 24722
rect 12514 24670 12516 24722
rect 12460 24164 12516 24670
rect 12796 24724 12852 24734
rect 12796 24630 12852 24668
rect 12460 24098 12516 24108
rect 13020 24162 13076 26460
rect 13356 24836 13412 24846
rect 13356 24834 13524 24836
rect 13356 24782 13358 24834
rect 13410 24782 13524 24834
rect 13356 24780 13524 24782
rect 13356 24770 13412 24780
rect 13020 24110 13022 24162
rect 13074 24110 13076 24162
rect 13020 24098 13076 24110
rect 12236 23938 12628 23940
rect 12236 23886 12238 23938
rect 12290 23886 12628 23938
rect 12236 23884 12628 23886
rect 12236 23874 12292 23884
rect 11900 23762 11956 23772
rect 12572 23154 12628 23884
rect 12796 23938 12852 23950
rect 12796 23886 12798 23938
rect 12850 23886 12852 23938
rect 12684 23828 12740 23866
rect 12684 23762 12740 23772
rect 12572 23102 12574 23154
rect 12626 23102 12628 23154
rect 12572 23090 12628 23102
rect 12684 23604 12740 23614
rect 12684 23266 12740 23548
rect 12684 23214 12686 23266
rect 12738 23214 12740 23266
rect 12236 23044 12292 23054
rect 12236 22950 12292 22988
rect 12684 22932 12740 23214
rect 12460 22876 12740 22932
rect 12012 22484 12068 22494
rect 12460 22484 12516 22876
rect 11788 22482 12516 22484
rect 11788 22430 12014 22482
rect 12066 22430 12516 22482
rect 11788 22428 12516 22430
rect 12012 22418 12068 22428
rect 11676 22316 11956 22372
rect 11900 21924 11956 22316
rect 12572 22370 12628 22382
rect 12572 22318 12574 22370
rect 12626 22318 12628 22370
rect 11564 21586 11620 21644
rect 11564 21534 11566 21586
rect 11618 21534 11620 21586
rect 11564 21522 11620 21534
rect 11788 21868 11900 21924
rect 11004 20972 11284 21028
rect 10892 20916 10948 20926
rect 10892 20822 10948 20860
rect 10332 20750 10334 20802
rect 10386 20750 10388 20802
rect 10332 20738 10388 20750
rect 9436 20486 9492 20524
rect 9996 20468 10052 20478
rect 9996 20132 10052 20412
rect 10108 20132 10164 20142
rect 9212 20076 9940 20132
rect 9996 20130 10164 20132
rect 9996 20078 10110 20130
rect 10162 20078 10164 20130
rect 9996 20076 10164 20078
rect 8428 18732 8596 18788
rect 8764 20018 8820 20030
rect 8764 19966 8766 20018
rect 8818 19966 8820 20018
rect 8764 19908 8820 19966
rect 9772 19908 9828 19918
rect 8428 18452 8484 18732
rect 8764 18564 8820 19852
rect 9660 19906 9828 19908
rect 9660 19854 9774 19906
rect 9826 19854 9828 19906
rect 9660 19852 9828 19854
rect 9660 19684 9716 19852
rect 9772 19842 9828 19852
rect 8876 19012 8932 19022
rect 9212 19012 9268 19022
rect 8932 19010 9268 19012
rect 8932 18958 9214 19010
rect 9266 18958 9268 19010
rect 8932 18956 9268 18958
rect 8876 18918 8932 18956
rect 9212 18946 9268 18956
rect 9660 18676 9716 19628
rect 9772 19236 9828 19246
rect 9772 19142 9828 19180
rect 9660 18610 9716 18620
rect 8876 18564 8932 18574
rect 8764 18508 8876 18564
rect 8204 18396 8484 18452
rect 8092 18340 8148 18350
rect 7868 18338 8148 18340
rect 7868 18286 8094 18338
rect 8146 18286 8148 18338
rect 7868 18284 8148 18286
rect 7868 17668 7924 18284
rect 8092 18274 8148 18284
rect 8204 18226 8260 18396
rect 8204 18174 8206 18226
rect 8258 18174 8260 18226
rect 8204 18162 8260 18174
rect 8652 17892 8708 17902
rect 8092 17780 8148 17790
rect 8092 17778 8372 17780
rect 8092 17726 8094 17778
rect 8146 17726 8372 17778
rect 8092 17724 8372 17726
rect 8092 17714 8148 17724
rect 7196 17614 7198 17666
rect 7250 17614 7252 17666
rect 6748 17108 6804 17118
rect 6748 16994 6804 17052
rect 6748 16942 6750 16994
rect 6802 16942 6804 16994
rect 6748 16930 6804 16942
rect 6860 16996 6916 17006
rect 6860 16902 6916 16940
rect 6972 16772 7028 17276
rect 7084 16996 7140 17006
rect 7084 16902 7140 16940
rect 6860 16716 7028 16772
rect 7196 16882 7252 17614
rect 7756 17666 7924 17668
rect 7756 17614 7870 17666
rect 7922 17614 7924 17666
rect 7756 17612 7924 17614
rect 7420 17108 7476 17118
rect 7476 17052 7588 17108
rect 7420 17042 7476 17052
rect 7532 16994 7588 17052
rect 7532 16942 7534 16994
rect 7586 16942 7588 16994
rect 7532 16930 7588 16942
rect 7756 17106 7812 17612
rect 7868 17602 7924 17612
rect 8204 17554 8260 17566
rect 8204 17502 8206 17554
rect 8258 17502 8260 17554
rect 8204 17444 8260 17502
rect 8204 17378 8260 17388
rect 7756 17054 7758 17106
rect 7810 17054 7812 17106
rect 7196 16830 7198 16882
rect 7250 16830 7252 16882
rect 6188 15986 6356 15988
rect 6188 15934 6190 15986
rect 6242 15934 6356 15986
rect 6188 15932 6356 15934
rect 6188 15922 6244 15932
rect 6188 15540 6244 15550
rect 6188 15426 6244 15484
rect 6188 15374 6190 15426
rect 6242 15374 6244 15426
rect 6188 15362 6244 15374
rect 5852 14590 5854 14642
rect 5906 14590 5908 14642
rect 5852 14578 5908 14590
rect 6300 15314 6356 15932
rect 6412 15988 6468 15998
rect 6636 15988 6692 15998
rect 6412 15986 6692 15988
rect 6412 15934 6414 15986
rect 6466 15934 6638 15986
rect 6690 15934 6692 15986
rect 6412 15932 6692 15934
rect 6412 15922 6468 15932
rect 6636 15922 6692 15932
rect 6748 15874 6804 15886
rect 6748 15822 6750 15874
rect 6802 15822 6804 15874
rect 6748 15428 6804 15822
rect 6860 15540 6916 16716
rect 6972 16100 7028 16110
rect 6972 16006 7028 16044
rect 7196 16098 7252 16830
rect 7196 16046 7198 16098
rect 7250 16046 7252 16098
rect 6860 15446 6916 15484
rect 7084 15988 7140 15998
rect 6748 15362 6804 15372
rect 6300 15262 6302 15314
rect 6354 15262 6356 15314
rect 6300 15204 6356 15262
rect 6300 14642 6356 15148
rect 6300 14590 6302 14642
rect 6354 14590 6356 14642
rect 6300 14578 6356 14590
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4956 11788 5460 11844
rect 5516 14532 5572 14542
rect 3052 10658 3108 10668
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 2044 5628 2772 5684
rect 2044 4562 2100 5628
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 2044 4510 2046 4562
rect 2098 4510 2100 4562
rect 2044 4498 2100 4510
rect 2492 4228 2548 4238
rect 2492 4134 2548 4172
rect 2940 4226 2996 4238
rect 2940 4174 2942 4226
rect 2994 4174 2996 4226
rect 2716 3666 2772 3678
rect 2716 3614 2718 3666
rect 2770 3614 2772 3666
rect 2044 3444 2100 3454
rect 1932 3442 2100 3444
rect 1932 3390 2046 3442
rect 2098 3390 2100 3442
rect 1932 3388 2100 3390
rect 2044 3378 2100 3388
rect 1708 2100 1764 3276
rect 1708 2034 1764 2044
rect 2716 800 2772 3614
rect 2940 3332 2996 4174
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4956 3554 5012 11788
rect 5516 9268 5572 14476
rect 6076 12066 6132 12078
rect 6076 12014 6078 12066
rect 6130 12014 6132 12066
rect 6076 11732 6132 12014
rect 6076 11666 6132 11676
rect 5516 9202 5572 9212
rect 7084 4338 7140 15932
rect 7196 15876 7252 16046
rect 7196 15810 7252 15820
rect 7420 16772 7476 16782
rect 7420 15538 7476 16716
rect 7756 16772 7812 17054
rect 7868 16884 7924 16894
rect 7868 16790 7924 16828
rect 7756 16706 7812 16716
rect 8204 16772 8260 16782
rect 7868 16100 7924 16110
rect 7868 16006 7924 16044
rect 8204 16098 8260 16716
rect 8204 16046 8206 16098
rect 8258 16046 8260 16098
rect 8204 16034 8260 16046
rect 8092 15988 8148 15998
rect 8092 15894 8148 15932
rect 7644 15876 7700 15886
rect 7700 15820 7812 15876
rect 7644 15782 7700 15820
rect 7420 15486 7422 15538
rect 7474 15486 7476 15538
rect 7420 15474 7476 15486
rect 7756 15540 7812 15820
rect 7756 15446 7812 15484
rect 8204 13636 8260 13646
rect 8204 12290 8260 13580
rect 8204 12238 8206 12290
rect 8258 12238 8260 12290
rect 8204 12226 8260 12238
rect 7084 4286 7086 4338
rect 7138 4286 7140 4338
rect 7084 4274 7140 4286
rect 5180 4116 5236 4126
rect 4956 3502 4958 3554
rect 5010 3502 5012 3554
rect 4956 3490 5012 3502
rect 5068 4114 5236 4116
rect 5068 4062 5182 4114
rect 5234 4062 5236 4114
rect 5068 4060 5236 4062
rect 5068 3332 5124 4060
rect 5180 4050 5236 4060
rect 2940 3266 2996 3276
rect 4732 3276 5124 3332
rect 6748 3666 6804 3678
rect 6748 3614 6750 3666
rect 6802 3614 6804 3666
rect 4732 800 4788 3276
rect 6748 800 6804 3614
rect 8316 3554 8372 17724
rect 8428 17556 8484 17566
rect 8428 17462 8484 17500
rect 8652 17554 8708 17836
rect 8652 17502 8654 17554
rect 8706 17502 8708 17554
rect 8652 17490 8708 17502
rect 8764 17554 8820 17566
rect 8764 17502 8766 17554
rect 8818 17502 8820 17554
rect 8540 17444 8596 17454
rect 8540 17106 8596 17388
rect 8540 17054 8542 17106
rect 8594 17054 8596 17106
rect 8540 17042 8596 17054
rect 8764 16772 8820 17502
rect 8764 16706 8820 16716
rect 8652 15988 8708 15998
rect 8652 15894 8708 15932
rect 8876 15148 8932 18508
rect 9772 18564 9828 18574
rect 9772 18470 9828 18508
rect 9772 18004 9828 18014
rect 9100 17892 9156 17902
rect 8988 17442 9044 17454
rect 8988 17390 8990 17442
rect 9042 17390 9044 17442
rect 8988 16996 9044 17390
rect 9100 17106 9156 17836
rect 9772 17780 9828 17948
rect 9212 17778 9828 17780
rect 9212 17726 9774 17778
rect 9826 17726 9828 17778
rect 9212 17724 9828 17726
rect 9212 17554 9268 17724
rect 9772 17714 9828 17724
rect 9212 17502 9214 17554
rect 9266 17502 9268 17554
rect 9212 17490 9268 17502
rect 9324 17554 9380 17566
rect 9324 17502 9326 17554
rect 9378 17502 9380 17554
rect 9100 17054 9102 17106
rect 9154 17054 9156 17106
rect 9100 17042 9156 17054
rect 8988 16930 9044 16940
rect 9324 16772 9380 17502
rect 9324 16706 9380 16716
rect 9772 16884 9828 16894
rect 9772 15988 9828 16828
rect 8428 15092 8932 15148
rect 9324 15986 9828 15988
rect 9324 15934 9774 15986
rect 9826 15934 9828 15986
rect 9324 15932 9828 15934
rect 8428 14196 8484 15092
rect 9324 14530 9380 15932
rect 9772 15922 9828 15932
rect 9884 15764 9940 20076
rect 10108 20066 10164 20076
rect 11004 20020 11060 20030
rect 10668 19908 10724 19918
rect 11004 19908 11060 19964
rect 10668 19814 10724 19852
rect 10892 19906 11060 19908
rect 10892 19854 11006 19906
rect 11058 19854 11060 19906
rect 10892 19852 11060 19854
rect 10668 19348 10724 19358
rect 10668 19254 10724 19292
rect 10108 19010 10164 19022
rect 10108 18958 10110 19010
rect 10162 18958 10164 19010
rect 10108 18564 10164 18958
rect 10108 18498 10164 18508
rect 10668 18564 10724 18574
rect 10892 18564 10948 19852
rect 11004 19842 11060 19852
rect 11004 19234 11060 19246
rect 11004 19182 11006 19234
rect 11058 19182 11060 19234
rect 11004 19012 11060 19182
rect 11004 18676 11060 18956
rect 11116 18676 11172 18686
rect 11004 18674 11172 18676
rect 11004 18622 11118 18674
rect 11170 18622 11172 18674
rect 11004 18620 11172 18622
rect 11116 18610 11172 18620
rect 10724 18508 10948 18564
rect 10668 18340 10724 18508
rect 10556 18338 10724 18340
rect 10556 18286 10670 18338
rect 10722 18286 10724 18338
rect 10556 18284 10724 18286
rect 10556 16324 10612 18284
rect 10668 18274 10724 18284
rect 11004 17332 11060 17342
rect 11004 17106 11060 17276
rect 11004 17054 11006 17106
rect 11058 17054 11060 17106
rect 11004 17042 11060 17054
rect 10556 16258 10612 16268
rect 10668 16994 10724 17006
rect 10668 16942 10670 16994
rect 10722 16942 10724 16994
rect 10668 16772 10724 16942
rect 9772 15708 9940 15764
rect 9996 16098 10052 16110
rect 9996 16046 9998 16098
rect 10050 16046 10052 16098
rect 9548 15540 9604 15550
rect 9548 15446 9604 15484
rect 9324 14478 9326 14530
rect 9378 14478 9380 14530
rect 9324 14466 9380 14478
rect 8988 14308 9044 14318
rect 9436 14308 9492 14318
rect 8988 14306 9492 14308
rect 8988 14254 8990 14306
rect 9042 14254 9438 14306
rect 9490 14254 9492 14306
rect 8988 14252 9492 14254
rect 8988 14242 9044 14252
rect 8428 14130 8484 14140
rect 9436 13412 9492 14252
rect 9660 14306 9716 14318
rect 9660 14254 9662 14306
rect 9714 14254 9716 14306
rect 9548 13860 9604 13870
rect 9660 13860 9716 14254
rect 9548 13858 9716 13860
rect 9548 13806 9550 13858
rect 9602 13806 9716 13858
rect 9548 13804 9716 13806
rect 9548 13794 9604 13804
rect 9660 13636 9716 13646
rect 9660 13542 9716 13580
rect 9772 13524 9828 15708
rect 9996 15540 10052 16046
rect 9996 15474 10052 15484
rect 10332 15426 10388 15438
rect 10332 15374 10334 15426
rect 10386 15374 10388 15426
rect 9884 15314 9940 15326
rect 9884 15262 9886 15314
rect 9938 15262 9940 15314
rect 9884 14196 9940 15262
rect 10108 15314 10164 15326
rect 10108 15262 10110 15314
rect 10162 15262 10164 15314
rect 10108 15148 10164 15262
rect 9884 14130 9940 14140
rect 9996 15092 10164 15148
rect 10332 15204 10388 15374
rect 10444 15428 10500 15438
rect 10668 15428 10724 16716
rect 10444 15426 10724 15428
rect 10444 15374 10446 15426
rect 10498 15374 10724 15426
rect 10444 15372 10724 15374
rect 10444 15362 10500 15372
rect 10332 15138 10388 15148
rect 10892 15204 10948 15242
rect 10892 15138 10948 15148
rect 9884 13860 9940 13870
rect 9996 13860 10052 15092
rect 11004 14532 11060 14542
rect 11228 14532 11284 20972
rect 11452 20578 11508 20590
rect 11452 20526 11454 20578
rect 11506 20526 11508 20578
rect 11340 19908 11396 19918
rect 11452 19908 11508 20526
rect 11676 20130 11732 20142
rect 11676 20078 11678 20130
rect 11730 20078 11732 20130
rect 11564 20020 11620 20030
rect 11676 20020 11732 20078
rect 11620 19964 11732 20020
rect 11564 19954 11620 19964
rect 11340 19906 11508 19908
rect 11340 19854 11342 19906
rect 11394 19854 11508 19906
rect 11340 19852 11508 19854
rect 11340 19572 11396 19852
rect 11340 19506 11396 19516
rect 11564 19460 11620 19470
rect 11788 19460 11844 21868
rect 11900 21858 11956 21868
rect 12012 22148 12068 22158
rect 12012 20914 12068 22092
rect 12236 21812 12292 21822
rect 12012 20862 12014 20914
rect 12066 20862 12068 20914
rect 12012 20850 12068 20862
rect 12124 21588 12180 21598
rect 11900 19908 11956 19918
rect 11900 19814 11956 19852
rect 11564 19458 11844 19460
rect 11564 19406 11566 19458
rect 11618 19406 11844 19458
rect 11564 19404 11844 19406
rect 11900 19572 11956 19582
rect 11564 19394 11620 19404
rect 11564 18564 11620 18574
rect 11564 18470 11620 18508
rect 11900 18450 11956 19516
rect 12012 19234 12068 19246
rect 12012 19182 12014 19234
rect 12066 19182 12068 19234
rect 12012 18564 12068 19182
rect 12124 19236 12180 21532
rect 12236 20242 12292 21756
rect 12572 21698 12628 22318
rect 12572 21646 12574 21698
rect 12626 21646 12628 21698
rect 12572 21252 12628 21646
rect 12572 21186 12628 21196
rect 12348 20916 12404 20926
rect 12348 20822 12404 20860
rect 12796 20916 12852 23886
rect 13468 21812 13524 24780
rect 13580 24164 13636 24174
rect 13580 23828 13636 24108
rect 13580 23268 13636 23772
rect 13580 22260 13636 23212
rect 13580 22166 13636 22204
rect 13468 21746 13524 21756
rect 13692 21476 13748 28252
rect 13804 23042 13860 28812
rect 13916 25396 13972 28924
rect 14028 28420 14084 28430
rect 14028 28082 14084 28364
rect 14028 28030 14030 28082
rect 14082 28030 14084 28082
rect 14028 27860 14084 28030
rect 14140 28082 14196 29036
rect 14252 28644 14308 29260
rect 14700 29314 14756 29326
rect 14700 29262 14702 29314
rect 14754 29262 14756 29314
rect 14588 28644 14644 28654
rect 14252 28642 14644 28644
rect 14252 28590 14590 28642
rect 14642 28590 14644 28642
rect 14252 28588 14644 28590
rect 14140 28030 14142 28082
rect 14194 28030 14196 28082
rect 14140 28018 14196 28030
rect 14252 27970 14308 27982
rect 14252 27918 14254 27970
rect 14306 27918 14308 27970
rect 14252 27860 14308 27918
rect 14028 27804 14308 27860
rect 14252 27076 14308 27086
rect 14476 27076 14532 27086
rect 14252 27074 14532 27076
rect 14252 27022 14254 27074
rect 14306 27022 14478 27074
rect 14530 27022 14532 27074
rect 14252 27020 14532 27022
rect 14252 26908 14308 27020
rect 14476 27010 14532 27020
rect 14588 26908 14644 28588
rect 14140 26852 14308 26908
rect 14364 26852 14420 26862
rect 14028 26292 14084 26302
rect 14028 25506 14084 26236
rect 14028 25454 14030 25506
rect 14082 25454 14084 25506
rect 14028 25442 14084 25454
rect 13916 24836 13972 25340
rect 13916 24770 13972 24780
rect 13916 23938 13972 23950
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13916 23604 13972 23886
rect 14028 23828 14084 23838
rect 14028 23734 14084 23772
rect 13916 23548 14084 23604
rect 14028 23268 14084 23548
rect 13804 22990 13806 23042
rect 13858 22990 13860 23042
rect 13804 22978 13860 22990
rect 13916 23212 14084 23268
rect 13804 22148 13860 22158
rect 13916 22148 13972 23212
rect 14028 23044 14084 23054
rect 14028 22372 14084 22988
rect 14028 22278 14084 22316
rect 13860 22092 13972 22148
rect 13804 22054 13860 22092
rect 13692 21420 13972 21476
rect 12908 21028 12964 21038
rect 12908 20934 12964 20972
rect 12796 20850 12852 20860
rect 12236 20190 12238 20242
rect 12290 20190 12292 20242
rect 12236 20178 12292 20190
rect 12572 20802 12628 20814
rect 12572 20750 12574 20802
rect 12626 20750 12628 20802
rect 12348 19684 12404 19694
rect 12348 19348 12404 19628
rect 12460 19460 12516 19470
rect 12572 19460 12628 20750
rect 13804 20578 13860 20590
rect 13804 20526 13806 20578
rect 13858 20526 13860 20578
rect 12908 20130 12964 20142
rect 12908 20078 12910 20130
rect 12962 20078 12964 20130
rect 12796 20018 12852 20030
rect 12796 19966 12798 20018
rect 12850 19966 12852 20018
rect 12796 19572 12852 19966
rect 12908 19908 12964 20078
rect 13804 20132 13860 20526
rect 12964 19852 13076 19908
rect 12908 19842 12964 19852
rect 12796 19506 12852 19516
rect 12460 19458 12572 19460
rect 12460 19406 12462 19458
rect 12514 19406 12572 19458
rect 12460 19404 12572 19406
rect 12460 19394 12516 19404
rect 12572 19366 12628 19404
rect 12348 19254 12404 19292
rect 13020 19348 13076 19852
rect 13804 19684 13860 20076
rect 13916 19684 13972 21420
rect 14140 21140 14196 26852
rect 14364 26758 14420 26796
rect 14476 26852 14644 26908
rect 14252 25396 14308 25406
rect 14252 25302 14308 25340
rect 14476 24276 14532 26852
rect 14700 26516 14756 29262
rect 14812 28866 14868 28878
rect 14812 28814 14814 28866
rect 14866 28814 14868 28866
rect 14812 27860 14868 28814
rect 15036 28644 15092 30156
rect 15148 30100 15204 30110
rect 15148 29538 15204 30044
rect 15148 29486 15150 29538
rect 15202 29486 15204 29538
rect 15148 29474 15204 29486
rect 15148 28644 15204 28654
rect 15036 28642 15204 28644
rect 15036 28590 15150 28642
rect 15202 28590 15204 28642
rect 15036 28588 15204 28590
rect 15148 28578 15204 28588
rect 14812 27766 14868 27804
rect 15036 28420 15092 28430
rect 15260 28420 15316 30268
rect 15484 30212 15540 32508
rect 15596 32498 15652 32508
rect 16044 31332 16100 31342
rect 16100 31276 16212 31332
rect 16044 31266 16100 31276
rect 15596 30996 15652 31006
rect 15596 30994 15876 30996
rect 15596 30942 15598 30994
rect 15650 30942 15876 30994
rect 15596 30940 15876 30942
rect 15596 30930 15652 30940
rect 15596 30212 15652 30222
rect 15484 30210 15652 30212
rect 15484 30158 15598 30210
rect 15650 30158 15652 30210
rect 15484 30156 15652 30158
rect 15484 28866 15540 30156
rect 15596 30146 15652 30156
rect 15708 30100 15764 30110
rect 15708 30006 15764 30044
rect 15820 29428 15876 30940
rect 16044 30882 16100 30894
rect 16044 30830 16046 30882
rect 16098 30830 16100 30882
rect 16044 30436 16100 30830
rect 16044 30370 16100 30380
rect 16156 30548 16212 31276
rect 15932 30212 15988 30222
rect 16156 30212 16212 30492
rect 15932 29538 15988 30156
rect 16044 30156 16212 30212
rect 16044 29652 16100 30156
rect 16268 29652 16324 38612
rect 16604 38162 16660 42588
rect 16940 42196 16996 42206
rect 16940 41972 16996 42140
rect 16828 41970 16996 41972
rect 16828 41918 16942 41970
rect 16994 41918 16996 41970
rect 16828 41916 16996 41918
rect 16828 41524 16884 41916
rect 16940 41906 16996 41916
rect 16828 41468 16996 41524
rect 16828 40516 16884 40526
rect 16828 39732 16884 40460
rect 16828 39638 16884 39676
rect 16716 39396 16772 39406
rect 16716 38946 16772 39340
rect 16716 38894 16718 38946
rect 16770 38894 16772 38946
rect 16716 38882 16772 38894
rect 16828 39058 16884 39070
rect 16828 39006 16830 39058
rect 16882 39006 16884 39058
rect 16828 38724 16884 39006
rect 16604 38110 16606 38162
rect 16658 38110 16660 38162
rect 16604 38098 16660 38110
rect 16716 38668 16884 38724
rect 16604 36932 16660 36942
rect 16604 36482 16660 36876
rect 16604 36430 16606 36482
rect 16658 36430 16660 36482
rect 16604 36418 16660 36430
rect 16380 36148 16436 36158
rect 16380 35922 16436 36092
rect 16380 35870 16382 35922
rect 16434 35870 16436 35922
rect 16380 35858 16436 35870
rect 16716 34132 16772 38668
rect 16716 34066 16772 34076
rect 16828 37154 16884 37166
rect 16828 37102 16830 37154
rect 16882 37102 16884 37154
rect 16828 35364 16884 37102
rect 16828 32676 16884 35308
rect 16940 32788 16996 41468
rect 17052 38612 17108 42812
rect 17276 42802 17332 42812
rect 17948 43314 18004 43326
rect 17948 43262 17950 43314
rect 18002 43262 18004 43314
rect 17836 42754 17892 42766
rect 17836 42702 17838 42754
rect 17890 42702 17892 42754
rect 17164 42644 17220 42654
rect 17836 42644 17892 42702
rect 17164 42642 17780 42644
rect 17164 42590 17166 42642
rect 17218 42590 17780 42642
rect 17164 42588 17780 42590
rect 17164 42578 17220 42588
rect 17388 42196 17444 42206
rect 17388 41970 17444 42140
rect 17724 42194 17780 42588
rect 17948 42644 18004 43262
rect 18060 42980 18116 43486
rect 18172 43316 18228 45612
rect 18172 43250 18228 43260
rect 18284 45444 18340 45454
rect 18060 42914 18116 42924
rect 18172 42754 18228 42766
rect 18172 42702 18174 42754
rect 18226 42702 18228 42754
rect 18172 42644 18228 42702
rect 17948 42588 18228 42644
rect 17836 42578 17892 42588
rect 17724 42142 17726 42194
rect 17778 42142 17780 42194
rect 17724 42130 17780 42142
rect 18172 42082 18228 42094
rect 18172 42030 18174 42082
rect 18226 42030 18228 42082
rect 17388 41918 17390 41970
rect 17442 41918 17444 41970
rect 17388 41906 17444 41918
rect 17724 41970 17780 41982
rect 17724 41918 17726 41970
rect 17778 41918 17780 41970
rect 17724 41188 17780 41918
rect 18060 41972 18116 41982
rect 18172 41972 18228 42030
rect 18060 41970 18228 41972
rect 18060 41918 18062 41970
rect 18114 41918 18228 41970
rect 18060 41916 18228 41918
rect 18060 41906 18116 41916
rect 17836 41188 17892 41198
rect 17724 41186 17892 41188
rect 17724 41134 17838 41186
rect 17890 41134 17892 41186
rect 17724 41132 17892 41134
rect 17836 41122 17892 41132
rect 18172 41076 18228 41086
rect 18172 40982 18228 41020
rect 17724 40962 17780 40974
rect 17724 40910 17726 40962
rect 17778 40910 17780 40962
rect 17724 40740 17780 40910
rect 18060 40962 18116 40974
rect 18060 40910 18062 40962
rect 18114 40910 18116 40962
rect 17780 40684 18004 40740
rect 17724 40674 17780 40684
rect 17388 39394 17444 39406
rect 17836 39396 17892 39406
rect 17388 39342 17390 39394
rect 17442 39342 17444 39394
rect 17388 39060 17444 39342
rect 17388 38994 17444 39004
rect 17500 39394 17892 39396
rect 17500 39342 17838 39394
rect 17890 39342 17892 39394
rect 17500 39340 17892 39342
rect 17500 38834 17556 39340
rect 17836 39330 17892 39340
rect 17500 38782 17502 38834
rect 17554 38782 17556 38834
rect 17500 38668 17556 38782
rect 17052 38546 17108 38556
rect 17388 38612 17556 38668
rect 17836 38836 17892 38846
rect 17836 38722 17892 38780
rect 17836 38670 17838 38722
rect 17890 38670 17892 38722
rect 17836 38658 17892 38670
rect 17164 36596 17220 36606
rect 17164 36482 17220 36540
rect 17164 36430 17166 36482
rect 17218 36430 17220 36482
rect 17164 36418 17220 36430
rect 17388 36482 17444 38612
rect 17612 38388 17668 38398
rect 17612 37378 17668 38332
rect 17612 37326 17614 37378
rect 17666 37326 17668 37378
rect 17612 37314 17668 37326
rect 17948 36596 18004 40684
rect 18060 40404 18116 40910
rect 18060 40338 18116 40348
rect 18060 39172 18116 39182
rect 18060 37380 18116 39116
rect 18284 38668 18340 45388
rect 18508 44212 18564 44222
rect 18396 44210 18564 44212
rect 18396 44158 18510 44210
rect 18562 44158 18564 44210
rect 18396 44156 18564 44158
rect 18396 42866 18452 44156
rect 18508 44146 18564 44156
rect 18396 42814 18398 42866
rect 18450 42814 18452 42866
rect 18396 42802 18452 42814
rect 18508 43652 18564 43662
rect 18508 43426 18564 43596
rect 18508 43374 18510 43426
rect 18562 43374 18564 43426
rect 18508 42644 18564 43374
rect 18732 43316 18788 43326
rect 18508 42578 18564 42588
rect 18620 42642 18676 42654
rect 18620 42590 18622 42642
rect 18674 42590 18676 42642
rect 18396 42532 18452 42542
rect 18396 42308 18452 42476
rect 18396 42252 18564 42308
rect 18508 42196 18564 42252
rect 18396 42084 18452 42094
rect 18396 41990 18452 42028
rect 18508 42082 18564 42140
rect 18508 42030 18510 42082
rect 18562 42030 18564 42082
rect 18508 42018 18564 42030
rect 18060 37286 18116 37324
rect 18172 38612 18340 38668
rect 18396 41860 18452 41870
rect 17388 36430 17390 36482
rect 17442 36430 17444 36482
rect 17388 35364 17444 36430
rect 17612 36540 18004 36596
rect 17500 35586 17556 35598
rect 17500 35534 17502 35586
rect 17554 35534 17556 35586
rect 17500 35476 17556 35534
rect 17500 35410 17556 35420
rect 17388 35298 17444 35308
rect 17612 33348 17668 36540
rect 17948 36370 18004 36382
rect 17948 36318 17950 36370
rect 18002 36318 18004 36370
rect 17948 36260 18004 36318
rect 17948 36194 18004 36204
rect 18060 35812 18116 35822
rect 18060 35586 18116 35756
rect 18172 35700 18228 38612
rect 18284 37042 18340 37054
rect 18284 36990 18286 37042
rect 18338 36990 18340 37042
rect 18284 36036 18340 36990
rect 18396 36482 18452 41804
rect 18620 41410 18676 42590
rect 18732 41860 18788 43260
rect 18844 42642 18900 42654
rect 18844 42590 18846 42642
rect 18898 42590 18900 42642
rect 18844 42308 18900 42590
rect 18844 42242 18900 42252
rect 18732 41794 18788 41804
rect 18844 42084 18900 42094
rect 18620 41358 18622 41410
rect 18674 41358 18676 41410
rect 18620 41346 18676 41358
rect 18508 41188 18564 41198
rect 18508 40628 18564 41132
rect 18732 41076 18788 41086
rect 18732 40982 18788 41020
rect 18620 40962 18676 40974
rect 18620 40910 18622 40962
rect 18674 40910 18676 40962
rect 18620 40740 18676 40910
rect 18620 40674 18676 40684
rect 18508 40562 18564 40572
rect 18844 39284 18900 42028
rect 18732 39228 18900 39284
rect 18620 38946 18676 38958
rect 18620 38894 18622 38946
rect 18674 38894 18676 38946
rect 18396 36430 18398 36482
rect 18450 36430 18452 36482
rect 18396 36418 18452 36430
rect 18508 38834 18564 38846
rect 18508 38782 18510 38834
rect 18562 38782 18564 38834
rect 18508 38724 18564 38782
rect 18620 38836 18676 38894
rect 18620 38770 18676 38780
rect 18732 38668 18788 39228
rect 18844 38948 18900 38958
rect 18844 38854 18900 38892
rect 18508 37044 18564 38668
rect 18620 38612 18788 38668
rect 18620 37490 18676 38612
rect 18620 37438 18622 37490
rect 18674 37438 18676 37490
rect 18620 37426 18676 37438
rect 18732 38050 18788 38062
rect 18732 37998 18734 38050
rect 18786 37998 18788 38050
rect 18732 37828 18788 37998
rect 18284 35980 18452 36036
rect 18284 35700 18340 35710
rect 18172 35698 18340 35700
rect 18172 35646 18286 35698
rect 18338 35646 18340 35698
rect 18172 35644 18340 35646
rect 18284 35634 18340 35644
rect 18060 35534 18062 35586
rect 18114 35534 18116 35586
rect 18060 35364 18116 35534
rect 18284 35476 18340 35486
rect 18396 35476 18452 35980
rect 18340 35420 18452 35476
rect 18284 35410 18340 35420
rect 18060 35298 18116 35308
rect 18508 35252 18564 36988
rect 18620 36148 18676 36158
rect 18620 35810 18676 36092
rect 18620 35758 18622 35810
rect 18674 35758 18676 35810
rect 18620 35476 18676 35758
rect 18620 35410 18676 35420
rect 18508 35196 18676 35252
rect 18620 34468 18676 35196
rect 18732 34914 18788 37772
rect 18844 37156 18900 37166
rect 18844 36260 18900 37100
rect 18956 36820 19012 45724
rect 19068 45666 19124 45678
rect 19068 45614 19070 45666
rect 19122 45614 19124 45666
rect 19068 45444 19124 45614
rect 20748 45666 20804 45678
rect 20748 45614 20750 45666
rect 20802 45614 20804 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19068 45378 19124 45388
rect 19180 44322 19236 44334
rect 19180 44270 19182 44322
rect 19234 44270 19236 44322
rect 19180 44100 19236 44270
rect 19740 44100 19796 44110
rect 19180 44098 19796 44100
rect 19180 44046 19742 44098
rect 19794 44046 19796 44098
rect 19180 44044 19796 44046
rect 19180 43652 19236 44044
rect 19740 44034 19796 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19180 43586 19236 43596
rect 19180 43426 19236 43438
rect 19180 43374 19182 43426
rect 19234 43374 19236 43426
rect 19180 42756 19236 43374
rect 20412 43428 20468 43438
rect 20412 43334 20468 43372
rect 19404 43316 19460 43326
rect 19404 43222 19460 43260
rect 19740 43314 19796 43326
rect 19740 43262 19742 43314
rect 19794 43262 19796 43314
rect 19740 42868 19796 43262
rect 20636 43314 20692 43326
rect 20636 43262 20638 43314
rect 20690 43262 20692 43314
rect 20636 43204 20692 43262
rect 20636 43138 20692 43148
rect 19740 42802 19796 42812
rect 19180 42700 19684 42756
rect 19404 42530 19460 42542
rect 19404 42478 19406 42530
rect 19458 42478 19460 42530
rect 19404 42308 19460 42478
rect 19404 42242 19460 42252
rect 19516 42532 19572 42542
rect 19516 42084 19572 42476
rect 19516 42018 19572 42028
rect 19628 42532 19684 42700
rect 19964 42532 20020 42542
rect 19628 42530 20020 42532
rect 19628 42478 19966 42530
rect 20018 42478 20020 42530
rect 19628 42476 20020 42478
rect 19404 41972 19460 41982
rect 19292 40962 19348 40974
rect 19292 40910 19294 40962
rect 19346 40910 19348 40962
rect 19292 40404 19348 40910
rect 19292 40338 19348 40348
rect 19180 38724 19236 38734
rect 19180 38630 19236 38668
rect 19404 38164 19460 41916
rect 19628 41860 19684 42476
rect 19964 42466 20020 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19404 38098 19460 38108
rect 19516 41804 19684 41860
rect 20076 42196 20132 42206
rect 19516 37268 19572 41804
rect 20076 41074 20132 42140
rect 20748 41972 20804 45614
rect 21532 45330 21588 46060
rect 21980 45890 22036 46060
rect 22876 46004 22932 49200
rect 22876 46002 23380 46004
rect 22876 45950 22878 46002
rect 22930 45950 23380 46002
rect 22876 45948 23380 45950
rect 22876 45938 22932 45948
rect 21980 45838 21982 45890
rect 22034 45838 22036 45890
rect 21980 45826 22036 45838
rect 23324 45890 23380 45948
rect 23324 45838 23326 45890
rect 23378 45838 23380 45890
rect 23324 45826 23380 45838
rect 24108 45892 24164 45902
rect 21756 45780 21812 45790
rect 21756 45666 21812 45724
rect 21756 45614 21758 45666
rect 21810 45614 21812 45666
rect 21756 45602 21812 45614
rect 23100 45668 23156 45678
rect 23100 45574 23156 45612
rect 21532 45278 21534 45330
rect 21586 45278 21588 45330
rect 21532 45266 21588 45278
rect 22764 44324 22820 44334
rect 20972 44212 21028 44222
rect 20972 43650 21028 44156
rect 22428 44212 22484 44222
rect 22428 44118 22484 44156
rect 22764 44210 22820 44268
rect 22764 44158 22766 44210
rect 22818 44158 22820 44210
rect 22764 44146 22820 44158
rect 23772 44212 23828 44222
rect 23772 44210 23940 44212
rect 23772 44158 23774 44210
rect 23826 44158 23940 44210
rect 23772 44156 23940 44158
rect 23772 44146 23828 44156
rect 21532 44098 21588 44110
rect 21532 44046 21534 44098
rect 21586 44046 21588 44098
rect 20972 43598 20974 43650
rect 21026 43598 21028 43650
rect 20972 43586 21028 43598
rect 21308 43652 21364 43662
rect 21308 43538 21364 43596
rect 21308 43486 21310 43538
rect 21362 43486 21364 43538
rect 21308 43474 21364 43486
rect 21532 43428 21588 44046
rect 21868 44098 21924 44110
rect 21868 44046 21870 44098
rect 21922 44046 21924 44098
rect 21868 43652 21924 44046
rect 21868 43586 21924 43596
rect 21420 43092 21476 43102
rect 21420 42866 21476 43036
rect 21420 42814 21422 42866
rect 21474 42814 21476 42866
rect 21420 42802 21476 42814
rect 20748 41906 20804 41916
rect 20076 41022 20078 41074
rect 20130 41022 20132 41074
rect 20076 41010 20132 41022
rect 20300 41186 20356 41198
rect 20300 41134 20302 41186
rect 20354 41134 20356 41186
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20300 39508 20356 41134
rect 20412 41076 20468 41086
rect 20412 40626 20468 41020
rect 20412 40574 20414 40626
rect 20466 40574 20468 40626
rect 20412 40562 20468 40574
rect 19628 39396 19684 39406
rect 19628 37490 19684 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20300 38948 20356 39452
rect 20636 40402 20692 40414
rect 20636 40350 20638 40402
rect 20690 40350 20692 40402
rect 20636 39396 20692 40350
rect 20636 39330 20692 39340
rect 21308 39396 21364 39406
rect 21308 39302 21364 39340
rect 20300 38882 20356 38892
rect 20300 37828 20356 37838
rect 20300 37734 20356 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37438 19630 37490
rect 19682 37438 19684 37490
rect 19628 37426 19684 37438
rect 20524 37380 20580 37390
rect 19516 37212 19684 37268
rect 19068 37156 19124 37166
rect 19068 37062 19124 37100
rect 19292 37044 19348 37054
rect 19292 36950 19348 36988
rect 18956 36764 19460 36820
rect 19404 36708 19460 36764
rect 19404 36652 19572 36708
rect 19292 36594 19348 36606
rect 19292 36542 19294 36594
rect 19346 36542 19348 36594
rect 19292 36484 19348 36542
rect 19348 36428 19460 36484
rect 19292 36418 19348 36428
rect 18844 35812 18900 36204
rect 19180 36372 19236 36382
rect 19180 35922 19236 36316
rect 19180 35870 19182 35922
rect 19234 35870 19236 35922
rect 19180 35858 19236 35870
rect 18844 35746 18900 35756
rect 19292 35812 19348 35822
rect 19292 35718 19348 35756
rect 18844 35588 18900 35598
rect 18900 35532 19012 35588
rect 18844 35494 18900 35532
rect 18732 34862 18734 34914
rect 18786 34862 18788 34914
rect 18732 34692 18788 34862
rect 18732 34626 18788 34636
rect 18620 34412 18788 34468
rect 18508 34356 18564 34366
rect 18172 34354 18564 34356
rect 18172 34302 18510 34354
rect 18562 34302 18564 34354
rect 18172 34300 18564 34302
rect 17724 33460 17780 33470
rect 17724 33366 17780 33404
rect 17500 33292 17668 33348
rect 17836 33348 17892 33358
rect 17052 33236 17108 33246
rect 17388 33236 17444 33246
rect 17108 33234 17444 33236
rect 17108 33182 17390 33234
rect 17442 33182 17444 33234
rect 17108 33180 17444 33182
rect 17052 33142 17108 33180
rect 17388 33170 17444 33180
rect 16940 32732 17220 32788
rect 16828 32620 16996 32676
rect 16716 30212 16772 30222
rect 16716 30118 16772 30156
rect 16604 30098 16660 30110
rect 16604 30046 16606 30098
rect 16658 30046 16660 30098
rect 16044 29558 16100 29596
rect 16156 29596 16324 29652
rect 16380 29764 16436 29774
rect 15932 29486 15934 29538
rect 15986 29486 15988 29538
rect 15932 29474 15988 29486
rect 15820 29362 15876 29372
rect 15484 28814 15486 28866
rect 15538 28814 15540 28866
rect 15484 28802 15540 28814
rect 15484 28644 15540 28654
rect 15484 28550 15540 28588
rect 15932 28420 15988 28430
rect 15260 28364 15652 28420
rect 15036 27858 15092 28364
rect 15036 27806 15038 27858
rect 15090 27806 15092 27858
rect 15036 26628 15092 27806
rect 15036 26572 15428 26628
rect 14700 26450 14756 26460
rect 14588 26292 14644 26302
rect 14588 24836 14644 26236
rect 15260 26292 15316 26302
rect 15260 26198 15316 26236
rect 14700 25956 14756 25966
rect 14700 25506 14756 25900
rect 14924 25620 14980 25630
rect 14924 25526 14980 25564
rect 14700 25454 14702 25506
rect 14754 25454 14756 25506
rect 14700 25442 14756 25454
rect 14812 25396 14868 25406
rect 14812 25302 14868 25340
rect 15036 25396 15092 25406
rect 15036 25302 15092 25340
rect 15148 25282 15204 25294
rect 15148 25230 15150 25282
rect 15202 25230 15204 25282
rect 15148 25172 15204 25230
rect 15260 25172 15316 25182
rect 15148 25116 15260 25172
rect 15260 25106 15316 25116
rect 14924 25060 14980 25070
rect 14812 24946 14868 24958
rect 14812 24894 14814 24946
rect 14866 24894 14868 24946
rect 14588 24780 14756 24836
rect 14364 24220 14532 24276
rect 14588 24610 14644 24622
rect 14588 24558 14590 24610
rect 14642 24558 14644 24610
rect 14364 23156 14420 24220
rect 14588 23828 14644 24558
rect 14588 23604 14644 23772
rect 14588 23538 14644 23548
rect 14700 23380 14756 24780
rect 14812 24612 14868 24894
rect 14812 24546 14868 24556
rect 14588 23324 14756 23380
rect 14364 23100 14532 23156
rect 14364 22484 14420 22494
rect 14364 22390 14420 22428
rect 14252 22260 14308 22270
rect 14252 22258 14420 22260
rect 14252 22206 14254 22258
rect 14306 22206 14420 22258
rect 14252 22204 14420 22206
rect 14252 22194 14308 22204
rect 14140 21074 14196 21084
rect 14364 20804 14420 22204
rect 14476 21588 14532 23100
rect 14476 21522 14532 21532
rect 14364 20710 14420 20748
rect 14588 21028 14644 23324
rect 14700 23154 14756 23166
rect 14700 23102 14702 23154
rect 14754 23102 14756 23154
rect 14700 22148 14756 23102
rect 14700 22082 14756 22092
rect 14924 21924 14980 25004
rect 15260 23268 15316 23278
rect 15260 23174 15316 23212
rect 15260 22820 15316 22830
rect 14364 20468 14420 20478
rect 13916 19628 14196 19684
rect 13804 19618 13860 19628
rect 14028 19460 14084 19470
rect 14028 19366 14084 19404
rect 12124 19142 12180 19180
rect 12012 18498 12068 18508
rect 13020 18562 13076 19292
rect 13804 19348 13860 19358
rect 13804 19254 13860 19292
rect 13020 18510 13022 18562
rect 13074 18510 13076 18562
rect 13020 18498 13076 18510
rect 13916 19236 13972 19246
rect 11900 18398 11902 18450
rect 11954 18398 11956 18450
rect 11900 18386 11956 18398
rect 13916 18450 13972 19180
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13916 18386 13972 18398
rect 13804 17332 13860 17342
rect 11788 17220 11844 17230
rect 11788 15316 11844 17164
rect 12908 16100 12964 16110
rect 12908 16006 12964 16044
rect 13244 16100 13300 16110
rect 13132 15876 13188 15886
rect 11788 15250 11844 15260
rect 12460 15652 12516 15662
rect 12460 15538 12516 15596
rect 12460 15486 12462 15538
rect 12514 15486 12516 15538
rect 12460 15148 12516 15486
rect 12796 15540 12852 15550
rect 12796 15446 12852 15484
rect 13132 15428 13188 15820
rect 13244 15538 13300 16044
rect 13804 16098 13860 17276
rect 13804 16046 13806 16098
rect 13858 16046 13860 16098
rect 13804 16034 13860 16046
rect 14028 16884 14084 16894
rect 14028 16212 14084 16828
rect 13468 15876 13524 15886
rect 13468 15782 13524 15820
rect 13244 15486 13246 15538
rect 13298 15486 13300 15538
rect 13244 15474 13300 15486
rect 12348 15092 12516 15148
rect 12908 15426 13188 15428
rect 12908 15374 13134 15426
rect 13186 15374 13188 15426
rect 12908 15372 13188 15374
rect 12908 15092 12964 15372
rect 13132 15362 13188 15372
rect 14028 15314 14084 16156
rect 14028 15262 14030 15314
rect 14082 15262 14084 15314
rect 14028 15250 14084 15262
rect 12012 14644 12068 14654
rect 12012 14550 12068 14588
rect 11004 14530 11508 14532
rect 11004 14478 11006 14530
rect 11058 14478 11508 14530
rect 11004 14476 11508 14478
rect 11004 14466 11060 14476
rect 11228 14306 11284 14318
rect 11228 14254 11230 14306
rect 11282 14254 11284 14306
rect 10780 14196 10836 14206
rect 9884 13858 10052 13860
rect 9884 13806 9886 13858
rect 9938 13806 10052 13858
rect 9884 13804 10052 13806
rect 10444 13858 10500 13870
rect 10444 13806 10446 13858
rect 10498 13806 10500 13858
rect 9884 13794 9940 13804
rect 10108 13748 10164 13758
rect 10444 13748 10500 13806
rect 10780 13858 10836 14140
rect 11228 14196 11284 14254
rect 11228 14130 11284 14140
rect 11452 13970 11508 14476
rect 12236 14308 12292 14318
rect 11452 13918 11454 13970
rect 11506 13918 11508 13970
rect 11452 13906 11508 13918
rect 12124 14306 12292 14308
rect 12124 14254 12238 14306
rect 12290 14254 12292 14306
rect 12124 14252 12292 14254
rect 10780 13806 10782 13858
rect 10834 13806 10836 13858
rect 10780 13794 10836 13806
rect 10108 13746 10500 13748
rect 10108 13694 10110 13746
rect 10162 13694 10500 13746
rect 10108 13692 10500 13694
rect 10108 13682 10164 13692
rect 9772 13468 9940 13524
rect 9436 13356 9828 13412
rect 8988 12178 9044 12190
rect 8988 12126 8990 12178
rect 9042 12126 9044 12178
rect 8988 12068 9044 12126
rect 9660 12068 9716 12078
rect 8988 12066 9716 12068
rect 8988 12014 9662 12066
rect 9714 12014 9716 12066
rect 8988 12012 9716 12014
rect 9436 11172 9492 11182
rect 9436 9938 9492 11116
rect 9436 9886 9438 9938
rect 9490 9886 9492 9938
rect 9436 9874 9492 9886
rect 8764 9828 8820 9838
rect 8764 9734 8820 9772
rect 9660 9828 9716 12012
rect 9772 11732 9828 13356
rect 9772 11666 9828 11676
rect 9660 9268 9716 9772
rect 9884 9716 9940 13468
rect 10444 12964 10500 13692
rect 12124 13636 12180 14252
rect 12236 14242 12292 14252
rect 12348 13860 12404 15092
rect 12572 15036 12964 15092
rect 13244 15090 13300 15102
rect 13244 15038 13246 15090
rect 13298 15038 13300 15090
rect 12460 14644 12516 14654
rect 12460 14418 12516 14588
rect 12572 14530 12628 15036
rect 12572 14478 12574 14530
rect 12626 14478 12628 14530
rect 12572 14466 12628 14478
rect 12460 14366 12462 14418
rect 12514 14366 12516 14418
rect 12460 14354 12516 14366
rect 11676 13580 12180 13636
rect 12236 13804 12740 13860
rect 10444 12898 10500 12908
rect 11452 12964 11508 12974
rect 11452 12292 11508 12908
rect 11676 12962 11732 13580
rect 11676 12910 11678 12962
rect 11730 12910 11732 12962
rect 11676 12898 11732 12910
rect 11900 12850 11956 12862
rect 11900 12798 11902 12850
rect 11954 12798 11956 12850
rect 11788 12738 11844 12750
rect 11788 12686 11790 12738
rect 11842 12686 11844 12738
rect 11452 12226 11508 12236
rect 11676 12404 11732 12414
rect 11564 11620 11620 11630
rect 11564 10498 11620 11564
rect 11564 10446 11566 10498
rect 11618 10446 11620 10498
rect 11564 10434 11620 10446
rect 11564 9940 11620 9950
rect 11676 9940 11732 12348
rect 11788 11172 11844 12686
rect 11900 12402 11956 12798
rect 11900 12350 11902 12402
rect 11954 12350 11956 12402
rect 11900 12338 11956 12350
rect 12124 12404 12180 12414
rect 12124 12310 12180 12348
rect 12236 12290 12292 13804
rect 12684 12964 12740 13804
rect 13244 13188 13300 15038
rect 13916 14308 13972 14318
rect 13916 14214 13972 14252
rect 14028 14306 14084 14318
rect 14028 14254 14030 14306
rect 14082 14254 14084 14306
rect 14028 13300 14084 14254
rect 14140 14084 14196 19628
rect 14364 19458 14420 20412
rect 14588 20468 14644 20972
rect 14588 20402 14644 20412
rect 14700 21868 14980 21924
rect 15148 22258 15204 22270
rect 15148 22206 15150 22258
rect 15202 22206 15204 22258
rect 14700 20130 14756 21868
rect 15148 21812 15204 22206
rect 15148 21746 15204 21756
rect 14924 21474 14980 21486
rect 14924 21422 14926 21474
rect 14978 21422 14980 21474
rect 14924 21252 14980 21422
rect 14924 21186 14980 21196
rect 14700 20078 14702 20130
rect 14754 20078 14756 20130
rect 14700 20066 14756 20078
rect 15148 20468 15204 20478
rect 14364 19406 14366 19458
rect 14418 19406 14420 19458
rect 14364 19394 14420 19406
rect 15148 19122 15204 20412
rect 15260 19908 15316 22764
rect 15372 22260 15428 26572
rect 15484 25172 15540 25182
rect 15484 24836 15540 25116
rect 15484 23714 15540 24780
rect 15484 23662 15486 23714
rect 15538 23662 15540 23714
rect 15484 23650 15540 23662
rect 15596 22484 15652 28364
rect 15932 28326 15988 28364
rect 16156 28196 16212 29596
rect 16268 29426 16324 29438
rect 16268 29374 16270 29426
rect 16322 29374 16324 29426
rect 16268 28756 16324 29374
rect 16268 28690 16324 28700
rect 16380 28644 16436 29708
rect 16380 28196 16436 28588
rect 15708 28140 16212 28196
rect 16268 28140 16436 28196
rect 16492 29316 16548 29326
rect 15708 25618 15764 28140
rect 16268 28084 16324 28140
rect 16156 28028 16324 28084
rect 15820 27858 15876 27870
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 15820 27300 15876 27806
rect 15820 27074 15876 27244
rect 15820 27022 15822 27074
rect 15874 27022 15876 27074
rect 15820 26290 15876 27022
rect 15820 26238 15822 26290
rect 15874 26238 15876 26290
rect 15820 26226 15876 26238
rect 15932 26962 15988 26974
rect 15932 26910 15934 26962
rect 15986 26910 15988 26962
rect 15708 25566 15710 25618
rect 15762 25566 15764 25618
rect 15708 25554 15764 25566
rect 15820 25844 15876 25854
rect 15708 25282 15764 25294
rect 15708 25230 15710 25282
rect 15762 25230 15764 25282
rect 15708 22596 15764 25230
rect 15820 22820 15876 25788
rect 15932 25732 15988 26910
rect 15932 25666 15988 25676
rect 16044 26404 16100 26414
rect 15932 25396 15988 25406
rect 15932 25302 15988 25340
rect 16044 24722 16100 26348
rect 16044 24670 16046 24722
rect 16098 24670 16100 24722
rect 16044 24658 16100 24670
rect 16156 24612 16212 28028
rect 16380 27972 16436 27982
rect 16380 27878 16436 27916
rect 16380 27074 16436 27086
rect 16380 27022 16382 27074
rect 16434 27022 16436 27074
rect 16380 26740 16436 27022
rect 16380 26674 16436 26684
rect 16268 26404 16324 26414
rect 16268 26310 16324 26348
rect 16492 25844 16548 29260
rect 16604 28644 16660 30046
rect 16716 29652 16772 29662
rect 16716 29558 16772 29596
rect 16828 28644 16884 28654
rect 16604 28642 16884 28644
rect 16604 28590 16830 28642
rect 16882 28590 16884 28642
rect 16604 28588 16884 28590
rect 16604 28420 16660 28430
rect 16604 28082 16660 28364
rect 16604 28030 16606 28082
rect 16658 28030 16660 28082
rect 16604 28018 16660 28030
rect 16828 27972 16884 28588
rect 16940 28196 16996 32620
rect 17052 28196 17108 28206
rect 16940 28140 17052 28196
rect 17052 28130 17108 28140
rect 16828 27906 16884 27916
rect 16716 27748 16772 27758
rect 16604 27188 16660 27198
rect 16604 26962 16660 27132
rect 16604 26910 16606 26962
rect 16658 26910 16660 26962
rect 16604 26898 16660 26910
rect 16716 26516 16772 27692
rect 17052 26962 17108 26974
rect 17052 26910 17054 26962
rect 17106 26910 17108 26962
rect 16940 26852 16996 26862
rect 16940 26758 16996 26796
rect 16716 26450 16772 26460
rect 16156 23268 16212 24556
rect 16268 25788 16548 25844
rect 16716 26180 16772 26190
rect 17052 26180 17108 26910
rect 16716 26178 17108 26180
rect 16716 26126 16718 26178
rect 16770 26126 17108 26178
rect 16716 26124 17108 26126
rect 16716 25844 16772 26124
rect 17164 26068 17220 32732
rect 17388 30884 17444 30894
rect 17388 29652 17444 30828
rect 17388 29586 17444 29596
rect 17388 28420 17444 28430
rect 17276 28364 17388 28420
rect 17276 26180 17332 28364
rect 17388 28326 17444 28364
rect 17276 26114 17332 26124
rect 17388 28196 17444 28206
rect 16268 23492 16324 25788
rect 16716 25778 16772 25788
rect 17052 26012 17220 26068
rect 16604 25732 16660 25742
rect 16492 25620 16548 25630
rect 16492 25526 16548 25564
rect 16492 25060 16548 25070
rect 16492 24946 16548 25004
rect 16492 24894 16494 24946
rect 16546 24894 16548 24946
rect 16492 24882 16548 24894
rect 16604 24946 16660 25676
rect 16604 24894 16606 24946
rect 16658 24894 16660 24946
rect 16604 24882 16660 24894
rect 16940 25732 16996 25742
rect 16380 24722 16436 24734
rect 16380 24670 16382 24722
rect 16434 24670 16436 24722
rect 16380 24612 16436 24670
rect 16380 24546 16436 24556
rect 16716 24724 16772 24734
rect 16604 24500 16660 24510
rect 16492 23828 16548 23838
rect 16492 23734 16548 23772
rect 16268 23436 16548 23492
rect 16156 23202 16212 23212
rect 15820 22754 15876 22764
rect 16380 23156 16436 23166
rect 15708 22530 15764 22540
rect 16380 22484 16436 23100
rect 15596 22418 15652 22428
rect 16268 22482 16436 22484
rect 16268 22430 16382 22482
rect 16434 22430 16436 22482
rect 16268 22428 16436 22430
rect 16044 22370 16100 22382
rect 16044 22318 16046 22370
rect 16098 22318 16100 22370
rect 15372 22204 15876 22260
rect 15372 22036 15428 22046
rect 15372 20802 15428 21980
rect 15708 21812 15764 21822
rect 15708 21698 15764 21756
rect 15708 21646 15710 21698
rect 15762 21646 15764 21698
rect 15708 21634 15764 21646
rect 15372 20750 15374 20802
rect 15426 20750 15428 20802
rect 15372 20738 15428 20750
rect 15596 21476 15652 21486
rect 15596 20916 15652 21420
rect 15596 20690 15652 20860
rect 15596 20638 15598 20690
rect 15650 20638 15652 20690
rect 15596 20626 15652 20638
rect 15372 20132 15428 20142
rect 15428 20076 15540 20132
rect 15372 20038 15428 20076
rect 15260 19852 15428 19908
rect 15260 19348 15316 19358
rect 15260 19234 15316 19292
rect 15260 19182 15262 19234
rect 15314 19182 15316 19234
rect 15260 19170 15316 19182
rect 15148 19070 15150 19122
rect 15202 19070 15204 19122
rect 15148 19058 15204 19070
rect 14924 19010 14980 19022
rect 14924 18958 14926 19010
rect 14978 18958 14980 19010
rect 14812 18340 14868 18350
rect 14364 16212 14420 16222
rect 14812 16212 14868 18284
rect 14364 16210 14868 16212
rect 14364 16158 14366 16210
rect 14418 16158 14868 16210
rect 14364 16156 14868 16158
rect 14364 16146 14420 16156
rect 14700 15986 14756 15998
rect 14700 15934 14702 15986
rect 14754 15934 14756 15986
rect 14252 15876 14308 15886
rect 14252 14532 14308 15820
rect 14700 15876 14756 15934
rect 14812 15986 14868 16156
rect 14812 15934 14814 15986
rect 14866 15934 14868 15986
rect 14812 15922 14868 15934
rect 14700 15810 14756 15820
rect 14924 15540 14980 18958
rect 15148 18676 15204 18686
rect 15148 18582 15204 18620
rect 15372 18452 15428 19852
rect 15484 18564 15540 20076
rect 15596 19012 15652 19022
rect 15596 19010 15764 19012
rect 15596 18958 15598 19010
rect 15650 18958 15764 19010
rect 15596 18956 15764 18958
rect 15596 18946 15652 18956
rect 15596 18564 15652 18574
rect 15484 18562 15652 18564
rect 15484 18510 15598 18562
rect 15650 18510 15652 18562
rect 15484 18508 15652 18510
rect 15596 18498 15652 18508
rect 15372 18396 15540 18452
rect 15036 17554 15092 17566
rect 15036 17502 15038 17554
rect 15090 17502 15092 17554
rect 15036 16884 15092 17502
rect 15036 16818 15092 16828
rect 15260 15986 15316 15998
rect 15260 15934 15262 15986
rect 15314 15934 15316 15986
rect 14924 15474 14980 15484
rect 15036 15874 15092 15886
rect 15036 15822 15038 15874
rect 15090 15822 15092 15874
rect 14588 15428 14644 15438
rect 14476 14980 14532 14990
rect 14364 14532 14420 14542
rect 14252 14530 14420 14532
rect 14252 14478 14366 14530
rect 14418 14478 14420 14530
rect 14252 14476 14420 14478
rect 14364 14466 14420 14476
rect 14252 14308 14308 14318
rect 14476 14308 14532 14924
rect 14588 14530 14644 15372
rect 14700 15202 14756 15214
rect 14700 15150 14702 15202
rect 14754 15150 14756 15202
rect 14700 15148 14756 15150
rect 14700 15092 14868 15148
rect 14812 14642 14868 15092
rect 14812 14590 14814 14642
rect 14866 14590 14868 14642
rect 14812 14578 14868 14590
rect 14588 14478 14590 14530
rect 14642 14478 14644 14530
rect 14588 14466 14644 14478
rect 15036 14530 15092 15822
rect 15260 15652 15316 15934
rect 15372 15988 15428 15998
rect 15372 15894 15428 15932
rect 15260 15586 15316 15596
rect 15036 14478 15038 14530
rect 15090 14478 15092 14530
rect 15036 14466 15092 14478
rect 15260 14420 15316 14430
rect 15260 14326 15316 14364
rect 14308 14252 14532 14308
rect 14252 14214 14308 14252
rect 14140 14028 14532 14084
rect 13804 13244 14084 13300
rect 13244 13132 13748 13188
rect 12684 12870 12740 12908
rect 13020 12964 13076 12974
rect 13356 12964 13412 12974
rect 13020 12962 13412 12964
rect 13020 12910 13022 12962
rect 13074 12910 13358 12962
rect 13410 12910 13412 12962
rect 13020 12908 13412 12910
rect 13020 12898 13076 12908
rect 13356 12898 13412 12908
rect 13692 12962 13748 13132
rect 13692 12910 13694 12962
rect 13746 12910 13748 12962
rect 13692 12898 13748 12910
rect 12460 12740 12516 12750
rect 12796 12740 12852 12750
rect 13580 12740 13636 12750
rect 12460 12738 12852 12740
rect 12460 12686 12462 12738
rect 12514 12686 12798 12738
rect 12850 12686 12852 12738
rect 12460 12684 12852 12686
rect 12460 12674 12516 12684
rect 12236 12238 12238 12290
rect 12290 12238 12292 12290
rect 12236 12226 12292 12238
rect 12796 11620 12852 12684
rect 13468 12738 13636 12740
rect 13468 12686 13582 12738
rect 13634 12686 13636 12738
rect 13468 12684 13636 12686
rect 13356 12292 13412 12302
rect 13356 12198 13412 12236
rect 13468 11620 13524 12684
rect 13580 12674 13636 12684
rect 13580 12292 13636 12302
rect 13804 12292 13860 13244
rect 13580 12290 13860 12292
rect 13580 12238 13582 12290
rect 13634 12238 13860 12290
rect 13580 12236 13860 12238
rect 13916 12962 13972 12974
rect 13916 12910 13918 12962
rect 13970 12910 13972 12962
rect 13916 12292 13972 12910
rect 14476 12850 14532 14028
rect 14588 12964 14644 12974
rect 14588 12870 14644 12908
rect 14476 12798 14478 12850
rect 14530 12798 14532 12850
rect 14252 12740 14308 12750
rect 13580 12226 13636 12236
rect 13916 12226 13972 12236
rect 14140 12738 14308 12740
rect 14140 12686 14254 12738
rect 14306 12686 14308 12738
rect 14140 12684 14308 12686
rect 14028 12180 14084 12190
rect 14140 12180 14196 12684
rect 14252 12674 14308 12684
rect 14476 12740 14532 12798
rect 14476 12684 14868 12740
rect 14028 12178 14196 12180
rect 14028 12126 14030 12178
rect 14082 12126 14196 12178
rect 14028 12124 14196 12126
rect 14028 12114 14084 12124
rect 13804 12066 13860 12078
rect 13804 12014 13806 12066
rect 13858 12014 13860 12066
rect 13468 11564 13748 11620
rect 12796 11554 12852 11564
rect 11788 11106 11844 11116
rect 13692 10722 13748 11564
rect 13692 10670 13694 10722
rect 13746 10670 13748 10722
rect 13692 10658 13748 10670
rect 13804 10500 13860 12014
rect 14476 11788 14532 12684
rect 14812 12402 14868 12684
rect 14812 12350 14814 12402
rect 14866 12350 14868 12402
rect 14812 12338 14868 12350
rect 13356 10444 13860 10500
rect 14364 11732 14532 11788
rect 15148 11732 15204 11742
rect 9884 9650 9940 9660
rect 11452 9938 11676 9940
rect 11452 9886 11566 9938
rect 11618 9886 11676 9938
rect 11452 9884 11676 9886
rect 9660 9202 9716 9212
rect 11452 9266 11508 9884
rect 11564 9874 11620 9884
rect 11676 9846 11732 9884
rect 12012 10388 12068 10398
rect 11452 9214 11454 9266
rect 11506 9214 11508 9266
rect 11452 9202 11508 9214
rect 11788 9268 11844 9278
rect 11788 9174 11844 9212
rect 12012 4338 12068 10332
rect 12460 10052 12516 10062
rect 12124 9940 12180 9950
rect 12124 9846 12180 9884
rect 12460 9826 12516 9996
rect 12460 9774 12462 9826
rect 12514 9774 12516 9826
rect 12348 9268 12404 9278
rect 12460 9268 12516 9774
rect 12348 9266 12516 9268
rect 12348 9214 12350 9266
rect 12402 9214 12516 9266
rect 12348 9212 12516 9214
rect 12572 9602 12628 9614
rect 12572 9550 12574 9602
rect 12626 9550 12628 9602
rect 12348 9202 12404 9212
rect 12012 4286 12014 4338
rect 12066 4286 12068 4338
rect 12012 4274 12068 4286
rect 8316 3502 8318 3554
rect 8370 3502 8372 3554
rect 8316 3490 8372 3502
rect 8764 4116 8820 4126
rect 8764 800 8820 4060
rect 9772 4116 9828 4126
rect 9772 4022 9828 4060
rect 12572 3554 12628 9550
rect 12684 9268 12740 9278
rect 12684 9042 12740 9212
rect 13356 9154 13412 10444
rect 14140 9940 14196 9950
rect 14140 9826 14196 9884
rect 14140 9774 14142 9826
rect 14194 9774 14196 9826
rect 14140 9762 14196 9774
rect 14364 9828 14420 11732
rect 14812 11620 14868 11630
rect 14812 11506 14868 11564
rect 14812 11454 14814 11506
rect 14866 11454 14868 11506
rect 14812 11442 14868 11454
rect 14924 10836 14980 10846
rect 15148 10836 15204 11676
rect 15484 11732 15540 18396
rect 15708 17332 15764 18956
rect 15708 17266 15764 17276
rect 15596 15874 15652 15886
rect 15596 15822 15598 15874
rect 15650 15822 15652 15874
rect 15596 15428 15652 15822
rect 15596 15362 15652 15372
rect 15484 11666 15540 11676
rect 15820 11620 15876 22204
rect 16044 21924 16100 22318
rect 16044 21364 16100 21868
rect 16044 21308 16212 21364
rect 16156 21252 16212 21308
rect 16156 21186 16212 21196
rect 16268 20804 16324 22428
rect 16380 22418 16436 22428
rect 16492 21812 16548 23436
rect 16604 22146 16660 24444
rect 16604 22094 16606 22146
rect 16658 22094 16660 22146
rect 16604 22082 16660 22094
rect 16716 22148 16772 24668
rect 16716 22082 16772 22092
rect 16604 21812 16660 21822
rect 16492 21810 16660 21812
rect 16492 21758 16606 21810
rect 16658 21758 16660 21810
rect 16492 21756 16660 21758
rect 16604 21746 16660 21756
rect 16716 21812 16772 21822
rect 16604 21586 16660 21598
rect 16604 21534 16606 21586
rect 16658 21534 16660 21586
rect 16268 20690 16324 20748
rect 16268 20638 16270 20690
rect 16322 20638 16324 20690
rect 16268 20626 16324 20638
rect 16380 21364 16436 21374
rect 16156 20468 16212 20478
rect 15932 20244 15988 20254
rect 15932 19458 15988 20188
rect 15932 19406 15934 19458
rect 15986 19406 15988 19458
rect 15932 19394 15988 19406
rect 16156 19346 16212 20412
rect 16156 19294 16158 19346
rect 16210 19294 16212 19346
rect 16156 19282 16212 19294
rect 16380 19348 16436 21308
rect 16604 21252 16660 21534
rect 16604 20018 16660 21196
rect 16604 19966 16606 20018
rect 16658 19966 16660 20018
rect 16604 19954 16660 19966
rect 16716 20244 16772 21756
rect 16268 18676 16324 18686
rect 16380 18676 16436 19292
rect 16716 19346 16772 20188
rect 16716 19294 16718 19346
rect 16770 19294 16772 19346
rect 16716 19282 16772 19294
rect 16268 18674 16436 18676
rect 16268 18622 16270 18674
rect 16322 18622 16436 18674
rect 16268 18620 16436 18622
rect 16268 18610 16324 18620
rect 16156 16660 16212 16670
rect 16156 16210 16212 16604
rect 16156 16158 16158 16210
rect 16210 16158 16212 16210
rect 16156 14532 16212 16158
rect 16940 15988 16996 25676
rect 17052 16772 17108 26012
rect 17388 25732 17444 28140
rect 17500 28084 17556 33292
rect 17836 33254 17892 33292
rect 17612 33122 17668 33134
rect 17612 33070 17614 33122
rect 17666 33070 17668 33122
rect 17612 32564 17668 33070
rect 17612 32498 17668 32508
rect 17948 33122 18004 33134
rect 17948 33070 17950 33122
rect 18002 33070 18004 33122
rect 17612 32340 17668 32350
rect 17612 32246 17668 32284
rect 17948 31108 18004 33070
rect 18172 32674 18228 34300
rect 18508 34290 18564 34300
rect 18172 32622 18174 32674
rect 18226 32622 18228 32674
rect 18172 32610 18228 32622
rect 18284 34132 18340 34142
rect 18620 34132 18676 34142
rect 18284 32674 18340 34076
rect 18508 34130 18676 34132
rect 18508 34078 18622 34130
rect 18674 34078 18676 34130
rect 18508 34076 18676 34078
rect 18508 34020 18564 34076
rect 18620 34066 18676 34076
rect 18508 33954 18564 33964
rect 18732 33908 18788 34412
rect 18956 34132 19012 35532
rect 19068 35586 19124 35598
rect 19068 35534 19070 35586
rect 19122 35534 19124 35586
rect 19068 34356 19124 35534
rect 19292 35476 19348 35486
rect 19180 34692 19236 34702
rect 19180 34598 19236 34636
rect 19068 34300 19236 34356
rect 19068 34132 19124 34142
rect 18956 34130 19124 34132
rect 18956 34078 19070 34130
rect 19122 34078 19124 34130
rect 18956 34076 19124 34078
rect 19068 34066 19124 34076
rect 18620 33852 18788 33908
rect 18844 34018 18900 34030
rect 18844 33966 18846 34018
rect 18898 33966 18900 34018
rect 18508 33348 18564 33358
rect 18508 33254 18564 33292
rect 18284 32622 18286 32674
rect 18338 32622 18340 32674
rect 18284 32610 18340 32622
rect 18060 32562 18116 32574
rect 18060 32510 18062 32562
rect 18114 32510 18116 32562
rect 18060 31780 18116 32510
rect 18060 31714 18116 31724
rect 18508 31668 18564 31678
rect 18172 31108 18228 31118
rect 17948 31052 18172 31108
rect 18172 31014 18228 31052
rect 18396 30994 18452 31006
rect 18396 30942 18398 30994
rect 18450 30942 18452 30994
rect 17836 30884 17892 30894
rect 18396 30884 18452 30942
rect 17836 30882 18452 30884
rect 17836 30830 17838 30882
rect 17890 30830 18452 30882
rect 17836 30828 18452 30830
rect 17612 29988 17668 29998
rect 17836 29988 17892 30828
rect 18508 30322 18564 31612
rect 18508 30270 18510 30322
rect 18562 30270 18564 30322
rect 18060 30212 18116 30222
rect 17612 29986 17836 29988
rect 17612 29934 17614 29986
rect 17666 29934 17836 29986
rect 17612 29932 17836 29934
rect 17612 29922 17668 29932
rect 17612 29316 17668 29326
rect 17612 29222 17668 29260
rect 17724 29092 17780 29932
rect 17836 29894 17892 29932
rect 17948 29986 18004 29998
rect 17948 29934 17950 29986
rect 18002 29934 18004 29986
rect 17948 29316 18004 29934
rect 17948 29250 18004 29260
rect 18060 29314 18116 30156
rect 18508 29988 18564 30270
rect 18396 29932 18564 29988
rect 18396 29428 18452 29932
rect 18508 29764 18564 29774
rect 18508 29650 18564 29708
rect 18508 29598 18510 29650
rect 18562 29598 18564 29650
rect 18508 29586 18564 29598
rect 18396 29372 18564 29428
rect 18060 29262 18062 29314
rect 18114 29262 18116 29314
rect 17724 29036 18004 29092
rect 17836 28642 17892 28654
rect 17836 28590 17838 28642
rect 17890 28590 17892 28642
rect 17836 28308 17892 28590
rect 17948 28420 18004 29036
rect 18060 28644 18116 29262
rect 18060 28578 18116 28588
rect 18172 28868 18228 28878
rect 17948 28364 18116 28420
rect 17836 28242 17892 28252
rect 17500 28028 17668 28084
rect 17500 27860 17556 27870
rect 17500 27766 17556 27804
rect 17500 27300 17556 27310
rect 17500 27074 17556 27244
rect 17500 27022 17502 27074
rect 17554 27022 17556 27074
rect 17500 27010 17556 27022
rect 17612 26908 17668 28028
rect 17948 27972 18004 27982
rect 17948 27878 18004 27916
rect 17276 25676 17444 25732
rect 17500 26852 17668 26908
rect 17164 25282 17220 25294
rect 17164 25230 17166 25282
rect 17218 25230 17220 25282
rect 17164 25060 17220 25230
rect 17164 23716 17220 25004
rect 17276 24500 17332 25676
rect 17276 24434 17332 24444
rect 17164 23650 17220 23660
rect 17388 23604 17444 23614
rect 17276 23380 17332 23390
rect 17276 20580 17332 23324
rect 17388 23266 17444 23548
rect 17500 23380 17556 26852
rect 17612 26740 17668 26750
rect 17612 26514 17668 26684
rect 17612 26462 17614 26514
rect 17666 26462 17668 26514
rect 17612 26450 17668 26462
rect 17724 25956 17780 25966
rect 17612 25732 17668 25742
rect 17612 25506 17668 25676
rect 17612 25454 17614 25506
rect 17666 25454 17668 25506
rect 17612 25442 17668 25454
rect 17724 25394 17780 25900
rect 17724 25342 17726 25394
rect 17778 25342 17780 25394
rect 17724 25330 17780 25342
rect 17836 25282 17892 25294
rect 17836 25230 17838 25282
rect 17890 25230 17892 25282
rect 17612 24948 17668 24958
rect 17612 24854 17668 24892
rect 17724 23938 17780 23950
rect 17724 23886 17726 23938
rect 17778 23886 17780 23938
rect 17500 23324 17668 23380
rect 17388 23214 17390 23266
rect 17442 23214 17444 23266
rect 17388 23202 17444 23214
rect 17500 23156 17556 23166
rect 17500 23062 17556 23100
rect 17276 20514 17332 20524
rect 17612 18564 17668 23324
rect 17724 23156 17780 23886
rect 17724 23090 17780 23100
rect 17612 18508 17780 18564
rect 17612 18340 17668 18350
rect 17612 18246 17668 18284
rect 17052 16210 17108 16716
rect 17500 16884 17556 16894
rect 17052 16158 17054 16210
rect 17106 16158 17108 16210
rect 17052 16146 17108 16158
rect 17388 16660 17444 16670
rect 17388 16098 17444 16604
rect 17388 16046 17390 16098
rect 17442 16046 17444 16098
rect 17388 16034 17444 16046
rect 16492 15874 16548 15886
rect 16492 15822 16494 15874
rect 16546 15822 16548 15874
rect 16156 14466 16212 14476
rect 16380 14532 16436 14542
rect 16268 14420 16324 14430
rect 16380 14420 16436 14476
rect 16268 14418 16436 14420
rect 16268 14366 16270 14418
rect 16322 14366 16436 14418
rect 16268 14364 16436 14366
rect 16268 14354 16324 14364
rect 15932 14306 15988 14318
rect 15932 14254 15934 14306
rect 15986 14254 15988 14306
rect 15932 14196 15988 14254
rect 15932 14130 15988 14140
rect 16492 14196 16548 15822
rect 16828 15204 16884 15214
rect 16940 15204 16996 15932
rect 17500 15538 17556 16828
rect 17724 16212 17780 18508
rect 17724 16146 17780 16156
rect 17500 15486 17502 15538
rect 17554 15486 17556 15538
rect 17500 15474 17556 15486
rect 16828 15202 16996 15204
rect 16828 15150 16830 15202
rect 16882 15150 16996 15202
rect 16828 15148 16996 15150
rect 16828 15138 16884 15148
rect 16492 14130 16548 14140
rect 17388 13076 17444 13086
rect 16716 12964 16772 12974
rect 16716 12870 16772 12908
rect 15596 11508 15652 11518
rect 15596 11394 15652 11452
rect 15596 11342 15598 11394
rect 15650 11342 15652 11394
rect 15596 11330 15652 11342
rect 15820 11394 15876 11564
rect 16492 11508 16548 11518
rect 16492 11414 16548 11452
rect 15820 11342 15822 11394
rect 15874 11342 15876 11394
rect 15820 11330 15876 11342
rect 16940 11396 16996 11406
rect 17388 11396 17444 13020
rect 16940 11394 17444 11396
rect 16940 11342 16942 11394
rect 16994 11342 17390 11394
rect 17442 11342 17444 11394
rect 16940 11340 17444 11342
rect 15932 11284 15988 11294
rect 15932 11282 16100 11284
rect 15932 11230 15934 11282
rect 15986 11230 16100 11282
rect 15932 11228 16100 11230
rect 15932 11218 15988 11228
rect 15820 10836 15876 10846
rect 14924 10834 15428 10836
rect 14924 10782 14926 10834
rect 14978 10782 15428 10834
rect 14924 10780 15428 10782
rect 14924 10770 14980 10780
rect 14364 9734 14420 9772
rect 14476 10610 14532 10622
rect 14476 10558 14478 10610
rect 14530 10558 14532 10610
rect 13356 9102 13358 9154
rect 13410 9102 13412 9154
rect 13356 9090 13412 9102
rect 13580 9714 13636 9726
rect 13580 9662 13582 9714
rect 13634 9662 13636 9714
rect 12684 8990 12686 9042
rect 12738 8990 12740 9042
rect 12684 8978 12740 8990
rect 13580 8428 13636 9662
rect 14476 9604 14532 10558
rect 15372 10610 15428 10780
rect 15372 10558 15374 10610
rect 15426 10558 15428 10610
rect 15372 10546 15428 10558
rect 15820 10610 15876 10780
rect 15820 10558 15822 10610
rect 15874 10558 15876 10610
rect 15820 10546 15876 10558
rect 15372 10388 15428 10398
rect 15372 10294 15428 10332
rect 15372 9940 15428 9950
rect 15372 9846 15428 9884
rect 15708 9828 15764 9838
rect 15484 9772 15708 9828
rect 14812 9604 14868 9614
rect 14476 9602 14868 9604
rect 14476 9550 14814 9602
rect 14866 9550 14868 9602
rect 14476 9548 14868 9550
rect 14812 9268 14868 9548
rect 14812 9202 14868 9212
rect 15484 8930 15540 9772
rect 15708 9734 15764 9772
rect 15932 9268 15988 9278
rect 15932 9174 15988 9212
rect 15484 8878 15486 8930
rect 15538 8878 15540 8930
rect 15484 8866 15540 8878
rect 13356 8372 13636 8428
rect 13356 4338 13412 8372
rect 13356 4286 13358 4338
rect 13410 4286 13412 4338
rect 13356 4274 13412 4286
rect 12572 3502 12574 3554
rect 12626 3502 12628 3554
rect 12572 3490 12628 3502
rect 12796 4116 12852 4126
rect 10780 3442 10836 3454
rect 10780 3390 10782 3442
rect 10834 3390 10836 3442
rect 10780 800 10836 3390
rect 12796 800 12852 4060
rect 14028 4116 14084 4126
rect 14028 4022 14084 4060
rect 16044 3554 16100 11228
rect 16492 10836 16548 10846
rect 16492 10742 16548 10780
rect 16940 9268 16996 11340
rect 17388 11330 17444 11340
rect 16828 9212 16940 9268
rect 16828 7698 16884 9212
rect 16940 9202 16996 9212
rect 17388 9716 17444 9726
rect 16828 7646 16830 7698
rect 16882 7646 16884 7698
rect 16828 6692 16884 7646
rect 17388 7362 17444 9660
rect 17388 7310 17390 7362
rect 17442 7310 17444 7362
rect 17388 7298 17444 7310
rect 16828 6626 16884 6636
rect 16044 3502 16046 3554
rect 16098 3502 16100 3554
rect 16044 3490 16100 3502
rect 17276 3666 17332 3678
rect 17276 3614 17278 3666
rect 17330 3614 17332 3666
rect 14812 3442 14868 3454
rect 14812 3390 14814 3442
rect 14866 3390 14868 3442
rect 14812 800 14868 3390
rect 17276 3388 17332 3614
rect 17836 3556 17892 25230
rect 17948 24948 18004 24958
rect 17948 24722 18004 24892
rect 17948 24670 17950 24722
rect 18002 24670 18004 24722
rect 17948 24658 18004 24670
rect 17948 23380 18004 23390
rect 18060 23380 18116 28364
rect 18172 28082 18228 28812
rect 18508 28420 18564 29372
rect 18508 28354 18564 28364
rect 18172 28030 18174 28082
rect 18226 28030 18228 28082
rect 18172 28018 18228 28030
rect 18508 28084 18564 28094
rect 18284 27972 18340 27982
rect 18172 27076 18228 27086
rect 18284 27076 18340 27916
rect 18396 27858 18452 27870
rect 18396 27806 18398 27858
rect 18450 27806 18452 27858
rect 18396 27300 18452 27806
rect 18396 27234 18452 27244
rect 18396 27076 18452 27086
rect 18284 27074 18452 27076
rect 18284 27022 18398 27074
rect 18450 27022 18452 27074
rect 18284 27020 18452 27022
rect 18172 26982 18228 27020
rect 18396 27010 18452 27020
rect 18508 26740 18564 28028
rect 18620 26964 18676 33852
rect 18844 31108 18900 33966
rect 18844 31042 18900 31052
rect 18956 33236 19012 33246
rect 18956 31218 19012 33180
rect 19180 32116 19236 34300
rect 19292 34242 19348 35420
rect 19292 34190 19294 34242
rect 19346 34190 19348 34242
rect 19292 34178 19348 34190
rect 19404 32788 19460 36428
rect 19516 34242 19572 36652
rect 19516 34190 19518 34242
rect 19570 34190 19572 34242
rect 19516 34178 19572 34190
rect 19628 33012 19684 37212
rect 20076 37154 20132 37166
rect 20076 37102 20078 37154
rect 20130 37102 20132 37154
rect 20076 37044 20132 37102
rect 20076 36978 20132 36988
rect 20524 37154 20580 37324
rect 20524 37102 20526 37154
rect 20578 37102 20580 37154
rect 20300 36932 20356 36942
rect 20300 36594 20356 36876
rect 20300 36542 20302 36594
rect 20354 36542 20356 36594
rect 20300 36530 20356 36542
rect 19852 36260 19908 36298
rect 19852 36194 19908 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19740 35812 19796 35822
rect 19740 35718 19796 35756
rect 20524 35028 20580 37102
rect 21420 37268 21476 37278
rect 20860 36596 20916 36606
rect 21420 36596 21476 37212
rect 20860 36502 20916 36540
rect 21196 36594 21476 36596
rect 21196 36542 21422 36594
rect 21474 36542 21476 36594
rect 21196 36540 21476 36542
rect 21196 36372 21252 36540
rect 21420 36530 21476 36540
rect 21196 35586 21252 36316
rect 21532 36260 21588 43372
rect 22092 43428 22148 43438
rect 22092 43426 22596 43428
rect 22092 43374 22094 43426
rect 22146 43374 22596 43426
rect 22092 43372 22596 43374
rect 22092 43362 22148 43372
rect 21868 43092 21924 43102
rect 21756 42642 21812 42654
rect 21756 42590 21758 42642
rect 21810 42590 21812 42642
rect 21756 42196 21812 42590
rect 21868 42642 21924 43036
rect 22540 42866 22596 43372
rect 22540 42814 22542 42866
rect 22594 42814 22596 42866
rect 22540 42802 22596 42814
rect 22652 42812 22932 42868
rect 22092 42756 22148 42766
rect 22316 42756 22372 42766
rect 22092 42754 22372 42756
rect 22092 42702 22094 42754
rect 22146 42702 22318 42754
rect 22370 42702 22372 42754
rect 22092 42700 22372 42702
rect 22092 42690 22148 42700
rect 22316 42690 22372 42700
rect 21868 42590 21870 42642
rect 21922 42590 21924 42642
rect 21868 42578 21924 42590
rect 22428 42308 22484 42318
rect 22316 42252 22428 42308
rect 21756 42130 21812 42140
rect 22204 42196 22260 42206
rect 22204 42082 22260 42140
rect 22316 42194 22372 42252
rect 22316 42142 22318 42194
rect 22370 42142 22372 42194
rect 22316 42130 22372 42142
rect 22204 42030 22206 42082
rect 22258 42030 22260 42082
rect 22204 42018 22260 42030
rect 22428 41748 22484 42252
rect 22652 42196 22708 42812
rect 22876 42754 22932 42812
rect 22876 42702 22878 42754
rect 22930 42702 22932 42754
rect 22876 42690 22932 42702
rect 23772 42754 23828 42766
rect 23772 42702 23774 42754
rect 23826 42702 23828 42754
rect 22764 42642 22820 42654
rect 22764 42590 22766 42642
rect 22818 42590 22820 42642
rect 22764 42196 22820 42590
rect 23436 42532 23492 42542
rect 23772 42532 23828 42702
rect 23436 42530 23828 42532
rect 23436 42478 23438 42530
rect 23490 42478 23828 42530
rect 23436 42476 23828 42478
rect 23884 42532 23940 44156
rect 24108 44210 24164 45836
rect 24220 44548 24276 49200
rect 25564 49140 25620 49200
rect 25900 49140 25956 49308
rect 25564 49084 25956 49140
rect 26236 46114 26292 49308
rect 26880 49200 26992 50000
rect 28224 49200 28336 50000
rect 29568 49200 29680 50000
rect 30912 49200 31024 50000
rect 32256 49200 32368 50000
rect 33600 49200 33712 50000
rect 34944 49200 35056 50000
rect 36288 49200 36400 50000
rect 37632 49200 37744 50000
rect 38976 49200 39088 50000
rect 40320 49200 40432 50000
rect 41664 49200 41776 50000
rect 43008 49200 43120 50000
rect 44352 49200 44464 50000
rect 45696 49200 45808 50000
rect 47040 49200 47152 50000
rect 26236 46062 26238 46114
rect 26290 46062 26292 46114
rect 26236 46050 26292 46062
rect 25228 45892 25284 45902
rect 25228 45798 25284 45836
rect 26908 45332 26964 49200
rect 28252 46116 28308 49200
rect 28252 46050 28308 46060
rect 29484 46116 29540 46126
rect 29484 46022 29540 46060
rect 28924 45892 28980 45902
rect 28924 45890 29204 45892
rect 28924 45838 28926 45890
rect 28978 45838 29204 45890
rect 28924 45836 29204 45838
rect 28924 45826 28980 45836
rect 26908 45266 26964 45276
rect 28140 45332 28196 45342
rect 28140 45238 28196 45276
rect 28476 45332 28532 45342
rect 25900 45220 25956 45230
rect 25900 45126 25956 45164
rect 24220 44482 24276 44492
rect 24332 45108 24388 45118
rect 24108 44158 24110 44210
rect 24162 44158 24164 44210
rect 24108 44146 24164 44158
rect 24220 43426 24276 43438
rect 24220 43374 24222 43426
rect 24274 43374 24276 43426
rect 23996 43092 24052 43102
rect 24220 43092 24276 43374
rect 24052 43036 24276 43092
rect 23996 42978 24052 43036
rect 23996 42926 23998 42978
rect 24050 42926 24052 42978
rect 23996 42914 24052 42926
rect 24332 42978 24388 45052
rect 25564 45108 25620 45118
rect 25564 45014 25620 45052
rect 27132 45108 27188 45118
rect 27132 45014 27188 45052
rect 25452 44548 25508 44558
rect 25452 44454 25508 44492
rect 28476 44546 28532 45276
rect 28476 44494 28478 44546
rect 28530 44494 28532 44546
rect 28476 44482 28532 44494
rect 27468 44436 27524 44446
rect 27468 44342 27524 44380
rect 27916 44436 27972 44446
rect 27916 44342 27972 44380
rect 24444 44324 24500 44334
rect 24444 44230 24500 44268
rect 28252 44322 28308 44334
rect 28252 44270 28254 44322
rect 28306 44270 28308 44322
rect 25340 43538 25396 43550
rect 25340 43486 25342 43538
rect 25394 43486 25396 43538
rect 24332 42926 24334 42978
rect 24386 42926 24388 42978
rect 24332 42914 24388 42926
rect 24780 43092 24836 43102
rect 24780 42866 24836 43036
rect 24780 42814 24782 42866
rect 24834 42814 24836 42866
rect 24780 42802 24836 42814
rect 23436 42466 23492 42476
rect 23436 42196 23492 42206
rect 22764 42140 23380 42196
rect 22652 42130 22708 42140
rect 22764 42028 23044 42084
rect 22540 41972 22596 41982
rect 22764 41972 22820 42028
rect 22540 41970 22820 41972
rect 22540 41918 22542 41970
rect 22594 41918 22820 41970
rect 22540 41916 22820 41918
rect 22988 41972 23044 42028
rect 23212 41972 23268 41982
rect 22988 41970 23268 41972
rect 22988 41918 23214 41970
rect 23266 41918 23268 41970
rect 22988 41916 23268 41918
rect 22540 41906 22596 41916
rect 23212 41906 23268 41916
rect 22876 41858 22932 41870
rect 22876 41806 22878 41858
rect 22930 41806 22932 41858
rect 22876 41748 22932 41806
rect 22428 41692 22932 41748
rect 22540 41076 22596 41086
rect 22540 40982 22596 41020
rect 22316 40964 22372 40974
rect 22316 40870 22372 40908
rect 22652 40964 22708 40974
rect 22652 40870 22708 40908
rect 22764 40740 22820 41692
rect 22876 41412 22932 41422
rect 22876 41186 22932 41356
rect 23212 41412 23268 41422
rect 23324 41412 23380 42140
rect 23436 41970 23492 42140
rect 23436 41918 23438 41970
rect 23490 41918 23492 41970
rect 23436 41906 23492 41918
rect 23548 41970 23604 41982
rect 23548 41918 23550 41970
rect 23602 41918 23604 41970
rect 23212 41410 23380 41412
rect 23212 41358 23214 41410
rect 23266 41358 23380 41410
rect 23212 41356 23380 41358
rect 23548 41412 23604 41918
rect 23212 41346 23268 41356
rect 23548 41346 23604 41356
rect 22876 41134 22878 41186
rect 22930 41134 22932 41186
rect 22876 41122 22932 41134
rect 22988 41300 23044 41310
rect 22988 40852 23044 41244
rect 23660 41188 23716 42476
rect 23884 42466 23940 42476
rect 23884 41970 23940 41982
rect 23884 41918 23886 41970
rect 23938 41918 23940 41970
rect 23884 41860 23940 41918
rect 23884 41794 23940 41804
rect 25340 41972 25396 43486
rect 26012 43426 26068 43438
rect 26012 43374 26014 43426
rect 26066 43374 26068 43426
rect 26012 42196 26068 43374
rect 26012 42130 26068 42140
rect 28140 43426 28196 43438
rect 28140 43374 28142 43426
rect 28194 43374 28196 43426
rect 28140 42084 28196 43374
rect 28252 43428 28308 44270
rect 29148 44210 29204 45836
rect 29596 44548 29652 49200
rect 30940 46116 30996 49200
rect 30940 46050 30996 46060
rect 32172 45892 32228 45902
rect 31836 45890 32228 45892
rect 31836 45838 32174 45890
rect 32226 45838 32228 45890
rect 31836 45836 32228 45838
rect 31836 45330 31892 45836
rect 32172 45826 32228 45836
rect 31836 45278 31838 45330
rect 31890 45278 31892 45330
rect 31836 45266 31892 45278
rect 31612 45108 31668 45118
rect 31612 45106 31780 45108
rect 31612 45054 31614 45106
rect 31666 45054 31780 45106
rect 31612 45052 31780 45054
rect 31612 45042 31668 45052
rect 30156 44996 30212 45006
rect 29596 44482 29652 44492
rect 30044 44994 30212 44996
rect 30044 44942 30158 44994
rect 30210 44942 30212 44994
rect 30044 44940 30212 44942
rect 29148 44158 29150 44210
rect 29202 44158 29204 44210
rect 29148 44146 29204 44158
rect 29372 44322 29428 44334
rect 29372 44270 29374 44322
rect 29426 44270 29428 44322
rect 28252 43362 28308 43372
rect 28700 43426 28756 43438
rect 28700 43374 28702 43426
rect 28754 43374 28756 43426
rect 28476 42756 28532 42766
rect 28476 42662 28532 42700
rect 28700 42084 28756 43374
rect 29036 43428 29092 43438
rect 28140 42018 28196 42028
rect 28476 42028 28756 42084
rect 28924 42980 28980 42990
rect 23772 41300 23828 41310
rect 23828 41244 24164 41300
rect 23772 41206 23828 41244
rect 23436 41132 23716 41188
rect 23100 41076 23156 41086
rect 23100 40982 23156 41020
rect 23212 40962 23268 40974
rect 23212 40910 23214 40962
rect 23266 40910 23268 40962
rect 23212 40852 23268 40910
rect 22988 40796 23268 40852
rect 23436 40740 23492 41132
rect 22652 40684 22820 40740
rect 23100 40684 23492 40740
rect 22092 40628 22148 40638
rect 21980 39508 22036 39518
rect 21980 39414 22036 39452
rect 21644 39396 21700 39406
rect 21644 39302 21700 39340
rect 21756 38722 21812 38734
rect 21756 38670 21758 38722
rect 21810 38670 21812 38722
rect 21756 37828 21812 38670
rect 21756 37762 21812 37772
rect 22092 37828 22148 40572
rect 22316 39620 22372 39630
rect 22316 39506 22372 39564
rect 22316 39454 22318 39506
rect 22370 39454 22372 39506
rect 22316 39442 22372 39454
rect 22428 39396 22484 39406
rect 22428 38050 22484 39340
rect 22428 37998 22430 38050
rect 22482 37998 22484 38050
rect 22428 37986 22484 37998
rect 22540 37828 22596 37838
rect 22092 37826 22596 37828
rect 22092 37774 22094 37826
rect 22146 37774 22542 37826
rect 22594 37774 22596 37826
rect 22092 37772 22596 37774
rect 22092 37762 22148 37772
rect 21196 35534 21198 35586
rect 21250 35534 21252 35586
rect 21196 35522 21252 35534
rect 21420 36258 21588 36260
rect 21420 36206 21534 36258
rect 21586 36206 21588 36258
rect 21420 36204 21588 36206
rect 20524 34972 21252 35028
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19964 34020 20020 34030
rect 19964 33926 20020 33964
rect 19628 32946 19684 32956
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19516 32788 19572 32798
rect 19404 32786 19908 32788
rect 19404 32734 19518 32786
rect 19570 32734 19908 32786
rect 19404 32732 19908 32734
rect 19516 32722 19572 32732
rect 19180 32060 19684 32116
rect 19404 31892 19460 31902
rect 19404 31798 19460 31836
rect 19068 31780 19124 31790
rect 19124 31724 19236 31780
rect 19068 31714 19124 31724
rect 18956 31166 18958 31218
rect 19010 31166 19012 31218
rect 18956 30100 19012 31166
rect 19068 31556 19124 31566
rect 19068 31218 19124 31500
rect 19068 31166 19070 31218
rect 19122 31166 19124 31218
rect 19068 31154 19124 31166
rect 19180 31218 19236 31724
rect 19180 31166 19182 31218
rect 19234 31166 19236 31218
rect 19180 31154 19236 31166
rect 19404 31554 19460 31566
rect 19404 31502 19406 31554
rect 19458 31502 19460 31554
rect 19404 31108 19460 31502
rect 19516 31554 19572 31566
rect 19516 31502 19518 31554
rect 19570 31502 19572 31554
rect 19516 31220 19572 31502
rect 19516 31154 19572 31164
rect 19404 31042 19460 31052
rect 19292 30994 19348 31006
rect 19292 30942 19294 30994
rect 19346 30942 19348 30994
rect 19180 30324 19236 30334
rect 18956 30034 19012 30044
rect 19068 30268 19180 30324
rect 18956 29876 19012 29886
rect 18956 29316 19012 29820
rect 18956 29222 19012 29260
rect 19068 29204 19124 30268
rect 19180 30258 19236 30268
rect 19180 29988 19236 29998
rect 19180 29894 19236 29932
rect 19068 29148 19236 29204
rect 18620 26898 18676 26908
rect 18732 28980 18788 28990
rect 18508 26674 18564 26684
rect 18004 23324 18116 23380
rect 18172 26180 18228 26190
rect 18172 23380 18228 26124
rect 18732 25508 18788 28924
rect 18956 28644 19012 28654
rect 18844 28308 18900 28318
rect 18844 27858 18900 28252
rect 18844 27806 18846 27858
rect 18898 27806 18900 27858
rect 18844 27794 18900 27806
rect 18956 27636 19012 28588
rect 18844 27580 19012 27636
rect 18844 26908 18900 27580
rect 19180 26962 19236 29148
rect 19292 28980 19348 30942
rect 19516 30994 19572 31006
rect 19516 30942 19518 30994
rect 19570 30942 19572 30994
rect 19516 30436 19572 30942
rect 19628 30884 19684 32060
rect 19852 31892 19908 32732
rect 20300 32452 20356 32462
rect 20300 32450 20468 32452
rect 20300 32398 20302 32450
rect 20354 32398 20468 32450
rect 20300 32396 20468 32398
rect 20300 32386 20356 32396
rect 19852 31826 19908 31836
rect 19740 31780 19796 31790
rect 19740 31686 19796 31724
rect 19964 31780 20020 31790
rect 19964 31686 20020 31724
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20300 31332 20356 31342
rect 19836 31322 20100 31332
rect 20188 31276 20300 31332
rect 19964 31220 20020 31230
rect 20188 31220 20244 31276
rect 20300 31266 20356 31276
rect 19964 31218 20244 31220
rect 19964 31166 19966 31218
rect 20018 31166 20244 31218
rect 19964 31164 20244 31166
rect 20412 31220 20468 32396
rect 19964 31154 20020 31164
rect 20300 31108 20356 31118
rect 20300 31014 20356 31052
rect 19628 30828 19796 30884
rect 19516 30370 19572 30380
rect 19628 30660 19684 30670
rect 19404 29764 19460 29774
rect 19404 29650 19460 29708
rect 19404 29598 19406 29650
rect 19458 29598 19460 29650
rect 19404 29586 19460 29598
rect 19628 29652 19684 30604
rect 19740 30324 19796 30828
rect 19740 30230 19796 30268
rect 20412 30324 20468 31164
rect 20524 31554 20580 31566
rect 20524 31502 20526 31554
rect 20578 31502 20580 31554
rect 20524 30436 20580 31502
rect 20636 30996 20692 31006
rect 20636 30902 20692 30940
rect 20748 30994 20804 31006
rect 20748 30942 20750 30994
rect 20802 30942 20804 30994
rect 20524 30370 20580 30380
rect 20412 30258 20468 30268
rect 20636 30324 20692 30334
rect 20748 30324 20804 30942
rect 20636 30322 20804 30324
rect 20636 30270 20638 30322
rect 20690 30270 20804 30322
rect 20636 30268 20804 30270
rect 20188 30100 20244 30110
rect 20076 29988 20132 30026
rect 20076 29922 20132 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19628 29596 20020 29652
rect 19964 29538 20020 29596
rect 19964 29486 19966 29538
rect 20018 29486 20020 29538
rect 19964 29474 20020 29486
rect 19516 29426 19572 29438
rect 19516 29374 19518 29426
rect 19570 29374 19572 29426
rect 19516 29316 19572 29374
rect 19628 29428 19684 29438
rect 19628 29334 19684 29372
rect 19740 29426 19796 29438
rect 19740 29374 19742 29426
rect 19794 29374 19796 29426
rect 19740 29316 19796 29374
rect 20188 29316 20244 30044
rect 20636 30100 20692 30268
rect 20636 30034 20692 30044
rect 19740 29260 20244 29316
rect 20412 29316 20468 29326
rect 19516 29250 19572 29260
rect 20412 29222 20468 29260
rect 21084 29316 21140 29326
rect 19292 28914 19348 28924
rect 19404 29204 19460 29214
rect 19180 26910 19182 26962
rect 19234 26910 19236 26962
rect 18844 26852 19012 26908
rect 18956 26516 19012 26852
rect 19180 26852 19236 26910
rect 19180 26786 19236 26796
rect 19292 28420 19348 28430
rect 19292 27858 19348 28364
rect 19292 27806 19294 27858
rect 19346 27806 19348 27858
rect 19292 27188 19348 27806
rect 18956 26460 19236 26516
rect 18956 26292 19012 26302
rect 18732 25452 18900 25508
rect 18620 25396 18676 25406
rect 18676 25340 18788 25396
rect 18620 25330 18676 25340
rect 18396 25284 18452 25294
rect 18396 25190 18452 25228
rect 18508 25172 18564 25182
rect 18508 24946 18564 25116
rect 18508 24894 18510 24946
rect 18562 24894 18564 24946
rect 18508 24882 18564 24894
rect 18284 24722 18340 24734
rect 18284 24670 18286 24722
rect 18338 24670 18340 24722
rect 18284 24612 18340 24670
rect 18396 24722 18452 24734
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 18396 24612 18452 24670
rect 18620 24724 18676 24734
rect 18620 24630 18676 24668
rect 18508 24612 18564 24622
rect 18396 24556 18508 24612
rect 18284 24052 18340 24556
rect 18508 24546 18564 24556
rect 18284 23996 18564 24052
rect 17948 23314 18004 23324
rect 18172 23314 18228 23324
rect 17948 23156 18004 23166
rect 18172 23156 18228 23166
rect 18004 23154 18228 23156
rect 18004 23102 18174 23154
rect 18226 23102 18228 23154
rect 18004 23100 18228 23102
rect 17948 22260 18004 23100
rect 18172 23090 18228 23100
rect 18508 22930 18564 23996
rect 18508 22878 18510 22930
rect 18562 22878 18564 22930
rect 18508 22866 18564 22878
rect 18620 23154 18676 23166
rect 18620 23102 18622 23154
rect 18674 23102 18676 23154
rect 18620 22708 18676 23102
rect 18508 22652 18676 22708
rect 18284 22484 18340 22494
rect 17948 20802 18004 22204
rect 18172 22482 18340 22484
rect 18172 22430 18286 22482
rect 18338 22430 18340 22482
rect 18172 22428 18340 22430
rect 18060 22148 18116 22158
rect 18060 20914 18116 22092
rect 18060 20862 18062 20914
rect 18114 20862 18116 20914
rect 18060 20850 18116 20862
rect 17948 20750 17950 20802
rect 18002 20750 18004 20802
rect 17948 20738 18004 20750
rect 18060 20020 18116 20030
rect 17948 19964 18060 20020
rect 17948 18564 18004 19964
rect 18060 19954 18116 19964
rect 18172 19236 18228 22428
rect 18284 22418 18340 22428
rect 18396 22258 18452 22270
rect 18396 22206 18398 22258
rect 18450 22206 18452 22258
rect 18284 22148 18340 22158
rect 18396 22148 18452 22206
rect 18340 22092 18452 22148
rect 18284 22082 18340 22092
rect 18508 22036 18564 22652
rect 18620 22484 18676 22494
rect 18732 22484 18788 25340
rect 18844 24836 18900 25452
rect 18956 25506 19012 26236
rect 18956 25454 18958 25506
rect 19010 25454 19012 25506
rect 18956 25442 19012 25454
rect 18844 24770 18900 24780
rect 19068 25060 19124 25070
rect 18620 22482 18732 22484
rect 18620 22430 18622 22482
rect 18674 22430 18732 22482
rect 18620 22428 18732 22430
rect 18620 22418 18676 22428
rect 18732 22390 18788 22428
rect 18844 23380 18900 23390
rect 18396 21980 18564 22036
rect 18396 21476 18452 21980
rect 18396 21410 18452 21420
rect 18060 19180 18228 19236
rect 18060 18788 18116 19180
rect 18172 19012 18228 19022
rect 18172 19010 18340 19012
rect 18172 18958 18174 19010
rect 18226 18958 18340 19010
rect 18172 18956 18340 18958
rect 18172 18946 18228 18956
rect 18060 18732 18228 18788
rect 18060 18564 18116 18574
rect 17948 18562 18116 18564
rect 17948 18510 18062 18562
rect 18114 18510 18116 18562
rect 17948 18508 18116 18510
rect 17948 18340 18004 18508
rect 18060 18498 18116 18508
rect 18172 18564 18228 18732
rect 18172 18470 18228 18508
rect 18284 18452 18340 18956
rect 18620 18564 18676 18574
rect 18508 18452 18564 18462
rect 18284 18450 18564 18452
rect 18284 18398 18510 18450
rect 18562 18398 18564 18450
rect 18284 18396 18564 18398
rect 17948 18274 18004 18284
rect 18060 18228 18116 18238
rect 18060 18134 18116 18172
rect 18396 17780 18452 17790
rect 18396 17666 18452 17724
rect 18396 17614 18398 17666
rect 18450 17614 18452 17666
rect 18396 17602 18452 17614
rect 18508 16884 18564 18396
rect 18620 17106 18676 18508
rect 18620 17054 18622 17106
rect 18674 17054 18676 17106
rect 18620 17042 18676 17054
rect 18844 17108 18900 23324
rect 19068 21812 19124 25004
rect 19180 24836 19236 26460
rect 19292 25508 19348 27132
rect 19404 27300 19460 29148
rect 19404 27074 19460 27244
rect 19404 27022 19406 27074
rect 19458 27022 19460 27074
rect 19404 27010 19460 27022
rect 19628 29204 19684 29214
rect 19404 26516 19460 26526
rect 19628 26516 19684 29148
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19852 27972 19908 27982
rect 19852 27878 19908 27916
rect 20412 27972 20468 27982
rect 20412 27878 20468 27916
rect 20524 27860 20580 27870
rect 20748 27860 20804 27870
rect 20580 27858 20804 27860
rect 20580 27806 20750 27858
rect 20802 27806 20804 27858
rect 20580 27804 20804 27806
rect 20524 27794 20580 27804
rect 19964 27748 20020 27758
rect 19964 27300 20020 27692
rect 19964 27186 20020 27244
rect 19964 27134 19966 27186
rect 20018 27134 20020 27186
rect 19964 27122 20020 27134
rect 20524 27300 20580 27310
rect 20412 27076 20468 27086
rect 20412 26982 20468 27020
rect 20300 26852 20356 26862
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19404 26514 19684 26516
rect 19404 26462 19406 26514
rect 19458 26462 19684 26514
rect 19404 26460 19684 26462
rect 19404 26450 19460 26460
rect 19628 26402 19684 26460
rect 19628 26350 19630 26402
rect 19682 26350 19684 26402
rect 19628 26338 19684 26350
rect 19852 26514 19908 26526
rect 19852 26462 19854 26514
rect 19906 26462 19908 26514
rect 19852 26292 19908 26462
rect 19852 26226 19908 26236
rect 19964 26516 20020 26526
rect 19964 26290 20020 26460
rect 19964 26238 19966 26290
rect 20018 26238 20020 26290
rect 19964 26226 20020 26238
rect 20300 26516 20356 26796
rect 20188 26180 20244 26190
rect 19516 25508 19572 25518
rect 19292 25506 19572 25508
rect 19292 25454 19518 25506
rect 19570 25454 19572 25506
rect 19292 25452 19572 25454
rect 19516 25442 19572 25452
rect 19740 25394 19796 25406
rect 19740 25342 19742 25394
rect 19794 25342 19796 25394
rect 19740 25284 19796 25342
rect 19740 25218 19796 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19852 24836 19908 24846
rect 19180 24780 19348 24836
rect 19180 24612 19236 24622
rect 19180 23828 19236 24556
rect 19180 23762 19236 23772
rect 19068 21746 19124 21756
rect 19292 19124 19348 24780
rect 19852 24742 19908 24780
rect 20188 24612 20244 26124
rect 20300 25394 20356 26460
rect 20300 25342 20302 25394
rect 20354 25342 20356 25394
rect 20300 25330 20356 25342
rect 20412 25506 20468 25518
rect 20412 25454 20414 25506
rect 20466 25454 20468 25506
rect 20412 24948 20468 25454
rect 20412 24882 20468 24892
rect 20300 24612 20356 24622
rect 20188 24610 20356 24612
rect 20188 24558 20302 24610
rect 20354 24558 20356 24610
rect 20188 24556 20356 24558
rect 20300 24546 20356 24556
rect 20188 23828 20244 23838
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19404 22484 19460 22494
rect 19460 22428 19684 22484
rect 19404 22418 19460 22428
rect 19628 21810 19684 22428
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21758 19630 21810
rect 19682 21758 19684 21810
rect 19628 21746 19684 21758
rect 19852 21700 19908 21710
rect 19404 21588 19460 21598
rect 19852 21588 19908 21644
rect 19460 21532 19908 21588
rect 19964 21586 20020 21598
rect 19964 21534 19966 21586
rect 20018 21534 20020 21586
rect 19404 21494 19460 21532
rect 19964 20692 20020 21534
rect 19964 20626 20020 20636
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19964 19348 20020 19358
rect 19404 19346 20020 19348
rect 19404 19294 19966 19346
rect 20018 19294 20020 19346
rect 19404 19292 20020 19294
rect 19404 19124 19460 19292
rect 19964 19282 20020 19292
rect 19292 19122 19460 19124
rect 19292 19070 19406 19122
rect 19458 19070 19460 19122
rect 19292 19068 19460 19070
rect 19180 19010 19236 19022
rect 19180 18958 19182 19010
rect 19234 18958 19236 19010
rect 19180 17666 19236 18958
rect 19292 18338 19348 18350
rect 19292 18286 19294 18338
rect 19346 18286 19348 18338
rect 19292 17780 19348 18286
rect 19404 18340 19460 19068
rect 19516 19124 19572 19134
rect 19516 19122 19684 19124
rect 19516 19070 19518 19122
rect 19570 19070 19684 19122
rect 19516 19068 19684 19070
rect 19516 19058 19572 19068
rect 19404 18274 19460 18284
rect 19516 18228 19572 18238
rect 19404 17780 19460 17790
rect 19292 17778 19460 17780
rect 19292 17726 19406 17778
rect 19458 17726 19460 17778
rect 19292 17724 19460 17726
rect 19404 17714 19460 17724
rect 19180 17614 19182 17666
rect 19234 17614 19236 17666
rect 19180 17602 19236 17614
rect 19516 17666 19572 18172
rect 19516 17614 19518 17666
rect 19570 17614 19572 17666
rect 19516 17602 19572 17614
rect 18844 17042 18900 17052
rect 19068 17556 19124 17566
rect 18508 16818 18564 16828
rect 18956 16994 19012 17006
rect 18956 16942 18958 16994
rect 19010 16942 19012 16994
rect 17948 16212 18004 16222
rect 17948 15148 18004 16156
rect 18956 15988 19012 16942
rect 19068 16772 19124 17500
rect 19404 17108 19460 17118
rect 19404 17014 19460 17052
rect 19628 16996 19684 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 17666 19796 17678
rect 19740 17614 19742 17666
rect 19794 17614 19796 17666
rect 19740 17556 19796 17614
rect 19740 17490 19796 17500
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 19852 17014 19908 17052
rect 19740 16996 19796 17006
rect 19628 16994 19796 16996
rect 19628 16942 19742 16994
rect 19794 16942 19796 16994
rect 19628 16940 19796 16942
rect 19068 16212 19124 16716
rect 19740 16212 19796 16940
rect 20076 16996 20132 17006
rect 20076 16902 20132 16940
rect 20188 16324 20244 23772
rect 20412 23268 20468 23278
rect 20524 23268 20580 27244
rect 20412 23266 20580 23268
rect 20412 23214 20414 23266
rect 20466 23214 20580 23266
rect 20412 23212 20580 23214
rect 20412 23202 20468 23212
rect 20300 23154 20356 23166
rect 20300 23102 20302 23154
rect 20354 23102 20356 23154
rect 20300 23044 20356 23102
rect 20300 19460 20356 22988
rect 20524 21476 20580 21486
rect 20524 21382 20580 21420
rect 20636 21028 20692 27804
rect 20748 27794 20804 27804
rect 20748 26290 20804 26302
rect 20748 26238 20750 26290
rect 20802 26238 20804 26290
rect 20748 25508 20804 26238
rect 20748 25442 20804 25452
rect 20860 24948 20916 24958
rect 20860 23380 20916 24892
rect 20860 23314 20916 23324
rect 20748 23042 20804 23054
rect 20748 22990 20750 23042
rect 20802 22990 20804 23042
rect 20748 21924 20804 22990
rect 21084 23044 21140 29260
rect 21196 28196 21252 34972
rect 21420 28420 21476 36204
rect 21532 36194 21588 36204
rect 22204 36370 22260 36382
rect 22204 36318 22206 36370
rect 22258 36318 22260 36370
rect 22204 35924 22260 36318
rect 22316 36372 22372 36382
rect 22316 36278 22372 36316
rect 22204 35858 22260 35868
rect 21980 35588 22036 35598
rect 21868 35532 21980 35588
rect 21644 34916 21700 34926
rect 21644 34018 21700 34860
rect 21644 33966 21646 34018
rect 21698 33966 21700 34018
rect 21644 33954 21700 33966
rect 21756 31892 21812 31902
rect 21532 31220 21588 31230
rect 21532 30994 21588 31164
rect 21532 30942 21534 30994
rect 21586 30942 21588 30994
rect 21532 30930 21588 30942
rect 21756 30994 21812 31836
rect 21756 30942 21758 30994
rect 21810 30942 21812 30994
rect 21756 30930 21812 30942
rect 21644 30548 21700 30558
rect 21644 30322 21700 30492
rect 21644 30270 21646 30322
rect 21698 30270 21700 30322
rect 21644 30258 21700 30270
rect 21756 28420 21812 28430
rect 21420 28364 21756 28420
rect 21196 28140 21588 28196
rect 21308 27524 21364 27534
rect 21308 27300 21364 27468
rect 21308 27206 21364 27244
rect 21196 27076 21252 27086
rect 21196 26908 21252 27020
rect 21420 26962 21476 26974
rect 21420 26910 21422 26962
rect 21474 26910 21476 26962
rect 21196 26852 21364 26908
rect 21196 26290 21252 26302
rect 21196 26238 21198 26290
rect 21250 26238 21252 26290
rect 21196 26180 21252 26238
rect 21196 26114 21252 26124
rect 21308 23492 21364 26852
rect 21420 26292 21476 26910
rect 21532 26908 21588 28140
rect 21644 27076 21700 28364
rect 21756 28354 21812 28364
rect 21868 27186 21924 35532
rect 21980 35522 22036 35532
rect 22428 35476 22484 37772
rect 22540 37762 22596 37772
rect 22652 36596 22708 40684
rect 22764 39508 22820 39518
rect 22764 38050 22820 39452
rect 22764 37998 22766 38050
rect 22818 37998 22820 38050
rect 22764 37986 22820 37998
rect 22652 36530 22708 36540
rect 22540 36260 22596 36270
rect 22540 36166 22596 36204
rect 22876 36258 22932 36270
rect 22876 36206 22878 36258
rect 22930 36206 22932 36258
rect 22876 35924 22932 36206
rect 22876 35858 22932 35868
rect 22428 35420 22596 35476
rect 22428 34916 22484 34926
rect 22428 34822 22484 34860
rect 22316 34804 22372 34814
rect 21980 33684 22036 33694
rect 21980 27300 22036 33628
rect 22316 31106 22372 34748
rect 22316 31054 22318 31106
rect 22370 31054 22372 31106
rect 22316 31042 22372 31054
rect 22316 28420 22372 28430
rect 22316 28082 22372 28364
rect 22316 28030 22318 28082
rect 22370 28030 22372 28082
rect 22316 28018 22372 28030
rect 22316 27636 22372 27646
rect 22204 27634 22372 27636
rect 22204 27582 22318 27634
rect 22370 27582 22372 27634
rect 22204 27580 22372 27582
rect 21980 27244 22148 27300
rect 21868 27134 21870 27186
rect 21922 27134 21924 27186
rect 21868 27122 21924 27134
rect 21644 27010 21700 27020
rect 21980 27076 22036 27114
rect 21980 27010 22036 27020
rect 21756 26962 21812 26974
rect 21756 26910 21758 26962
rect 21810 26910 21812 26962
rect 21532 26852 21700 26908
rect 21532 26516 21588 26526
rect 21532 26402 21588 26460
rect 21532 26350 21534 26402
rect 21586 26350 21588 26402
rect 21532 26338 21588 26350
rect 21420 26226 21476 26236
rect 21644 25172 21700 26852
rect 21756 26628 21812 26910
rect 22092 26908 22148 27244
rect 21756 26562 21812 26572
rect 21868 26852 22148 26908
rect 21868 25956 21924 26852
rect 21980 26786 22036 26796
rect 21980 26292 22036 26302
rect 21980 26198 22036 26236
rect 21868 25890 21924 25900
rect 22092 26068 22148 26078
rect 21308 23426 21364 23436
rect 21420 25116 21700 25172
rect 21196 23154 21252 23166
rect 21196 23102 21198 23154
rect 21250 23102 21252 23154
rect 21196 23044 21252 23102
rect 21140 22988 21252 23044
rect 21084 22978 21140 22988
rect 20860 22148 20916 22158
rect 20860 22054 20916 22092
rect 21308 22148 21364 22158
rect 21308 22054 21364 22092
rect 20748 21858 20804 21868
rect 20748 21700 20804 21710
rect 20748 21606 20804 21644
rect 20524 20972 20692 21028
rect 21084 21586 21140 21598
rect 21308 21588 21364 21598
rect 21084 21534 21086 21586
rect 21138 21534 21140 21586
rect 21084 21476 21140 21534
rect 20412 20692 20468 20702
rect 20412 20598 20468 20636
rect 20412 19906 20468 19918
rect 20412 19854 20414 19906
rect 20466 19854 20468 19906
rect 20412 19684 20468 19854
rect 20412 19618 20468 19628
rect 20300 19404 20468 19460
rect 20300 17556 20356 17566
rect 20300 16994 20356 17500
rect 20300 16942 20302 16994
rect 20354 16942 20356 16994
rect 20300 16930 20356 16942
rect 20188 16258 20244 16268
rect 20076 16212 20132 16222
rect 19740 16156 20020 16212
rect 19068 16146 19124 16156
rect 19740 15988 19796 15998
rect 18956 15148 19012 15932
rect 19628 15932 19740 15988
rect 19964 15988 20020 16156
rect 20076 16118 20132 16156
rect 19964 15932 20356 15988
rect 19628 15428 19684 15932
rect 19740 15922 19796 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19852 15540 19908 15550
rect 20300 15540 20356 15932
rect 19852 15538 20132 15540
rect 19852 15486 19854 15538
rect 19906 15486 20132 15538
rect 19852 15484 20132 15486
rect 19852 15474 19908 15484
rect 19740 15428 19796 15438
rect 19628 15426 19796 15428
rect 19628 15374 19742 15426
rect 19794 15374 19796 15426
rect 19628 15372 19796 15374
rect 19740 15362 19796 15372
rect 19964 15316 20020 15326
rect 17948 15092 18340 15148
rect 18284 14644 18340 15092
rect 18844 15092 19012 15148
rect 19404 15204 19460 15242
rect 19404 15138 19460 15148
rect 18284 14642 18788 14644
rect 18284 14590 18286 14642
rect 18338 14590 18788 14642
rect 18284 14588 18788 14590
rect 18284 14578 18340 14588
rect 18732 14418 18788 14588
rect 18844 14530 18900 15092
rect 19852 15090 19908 15102
rect 19852 15038 19854 15090
rect 19906 15038 19908 15090
rect 19852 14756 19908 15038
rect 19852 14690 19908 14700
rect 19964 14754 20020 15260
rect 20076 15204 20132 15484
rect 20076 15138 20132 15148
rect 20188 15538 20356 15540
rect 20188 15486 20302 15538
rect 20354 15486 20356 15538
rect 20188 15484 20356 15486
rect 19964 14702 19966 14754
rect 20018 14702 20020 14754
rect 19964 14690 20020 14702
rect 20188 14644 20244 15484
rect 20300 15474 20356 15484
rect 20412 15148 20468 19404
rect 20524 16660 20580 20972
rect 21084 20356 21140 21420
rect 21084 20290 21140 20300
rect 21196 21586 21364 21588
rect 21196 21534 21310 21586
rect 21362 21534 21364 21586
rect 21196 21532 21364 21534
rect 20748 20018 20804 20030
rect 20748 19966 20750 20018
rect 20802 19966 20804 20018
rect 20748 19684 20804 19966
rect 20748 19618 20804 19628
rect 20748 17780 20804 17790
rect 20748 17686 20804 17724
rect 20860 17220 20916 17230
rect 20748 16996 20804 17006
rect 20748 16902 20804 16940
rect 20860 16994 20916 17164
rect 20860 16942 20862 16994
rect 20914 16942 20916 16994
rect 20860 16930 20916 16942
rect 20636 16882 20692 16894
rect 21084 16884 21140 16894
rect 20636 16830 20638 16882
rect 20690 16830 20692 16882
rect 20636 16772 20692 16830
rect 20972 16882 21140 16884
rect 20972 16830 21086 16882
rect 21138 16830 21140 16882
rect 20972 16828 21140 16830
rect 20972 16772 21028 16828
rect 21084 16818 21140 16828
rect 20636 16716 21028 16772
rect 20524 16604 20804 16660
rect 20076 14588 20244 14644
rect 20300 15092 20468 15148
rect 20636 15874 20692 15886
rect 20636 15822 20638 15874
rect 20690 15822 20692 15874
rect 20636 15538 20692 15822
rect 20636 15486 20638 15538
rect 20690 15486 20692 15538
rect 18844 14478 18846 14530
rect 18898 14478 18900 14530
rect 18844 14466 18900 14478
rect 19068 14532 19124 14542
rect 18732 14366 18734 14418
rect 18786 14366 18788 14418
rect 18732 14354 18788 14366
rect 18508 14308 18564 14318
rect 18508 14306 18676 14308
rect 18508 14254 18510 14306
rect 18562 14254 18676 14306
rect 18508 14252 18676 14254
rect 18508 14242 18564 14252
rect 18620 13300 18676 14252
rect 18620 13244 19012 13300
rect 18956 12290 19012 13244
rect 18956 12238 18958 12290
rect 19010 12238 19012 12290
rect 18956 12226 19012 12238
rect 18844 12178 18900 12190
rect 18844 12126 18846 12178
rect 18898 12126 18900 12178
rect 18060 12068 18116 12078
rect 18844 12068 18900 12126
rect 19068 12068 19124 14476
rect 19852 14532 19908 14542
rect 20076 14532 20132 14588
rect 19852 14530 20132 14532
rect 19852 14478 19854 14530
rect 19906 14478 20132 14530
rect 19852 14476 20132 14478
rect 19852 14466 19908 14476
rect 20076 14420 20132 14476
rect 20076 14354 20132 14364
rect 19628 14308 19684 14318
rect 19964 14308 20020 14346
rect 19628 14306 19964 14308
rect 19628 14254 19630 14306
rect 19682 14254 19964 14306
rect 19628 14252 19964 14254
rect 19628 14242 19684 14252
rect 19964 14242 20020 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20300 13860 20356 15092
rect 20412 14420 20468 14430
rect 20412 14362 20468 14364
rect 20412 14310 20414 14362
rect 20466 14310 20468 14362
rect 20412 14298 20468 14310
rect 20524 14306 20580 14318
rect 20188 13804 20356 13860
rect 20524 14254 20526 14306
rect 20578 14254 20580 14306
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19292 12178 19348 12190
rect 19292 12126 19294 12178
rect 19346 12126 19348 12178
rect 18844 12012 19124 12068
rect 19180 12068 19236 12078
rect 18060 11506 18116 12012
rect 19180 11974 19236 12012
rect 18060 11454 18062 11506
rect 18114 11454 18116 11506
rect 18060 11442 18116 11454
rect 19180 10836 19236 10846
rect 19292 10836 19348 12126
rect 20188 11506 20244 13804
rect 20524 13748 20580 14254
rect 20524 13682 20580 13692
rect 20300 13636 20356 13646
rect 20300 13076 20356 13580
rect 20300 12982 20356 13020
rect 20524 12292 20580 12302
rect 20188 11454 20190 11506
rect 20242 11454 20244 11506
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19180 10834 19348 10836
rect 19180 10782 19182 10834
rect 19234 10782 19348 10834
rect 19180 10780 19348 10782
rect 20076 10836 20132 10846
rect 20188 10836 20244 11454
rect 20076 10834 20244 10836
rect 20076 10782 20078 10834
rect 20130 10782 20244 10834
rect 20076 10780 20244 10782
rect 20300 12236 20524 12292
rect 19180 10770 19236 10780
rect 19404 10724 19460 10734
rect 19404 10630 19460 10668
rect 20076 10724 20132 10780
rect 20076 10658 20132 10668
rect 19516 10610 19572 10622
rect 19516 10558 19518 10610
rect 19570 10558 19572 10610
rect 19516 10164 19572 10558
rect 19516 10108 20132 10164
rect 19964 9940 20020 9950
rect 19292 9938 20020 9940
rect 19292 9886 19966 9938
rect 20018 9886 20020 9938
rect 19292 9884 20020 9886
rect 18620 9716 18676 9726
rect 18620 9266 18676 9660
rect 18620 9214 18622 9266
rect 18674 9214 18676 9266
rect 18620 9202 18676 9214
rect 19180 9042 19236 9054
rect 19180 8990 19182 9042
rect 19234 8990 19236 9042
rect 19180 8932 19236 8990
rect 19292 9042 19348 9884
rect 19964 9874 20020 9884
rect 20076 9828 20132 10108
rect 20300 10050 20356 12236
rect 20524 12198 20580 12236
rect 20636 12180 20692 15486
rect 20748 15148 20804 16604
rect 20860 15876 20916 15886
rect 21196 15876 21252 21532
rect 21308 21522 21364 21532
rect 21308 20020 21364 20030
rect 21308 19926 21364 19964
rect 21420 19124 21476 25116
rect 21532 23268 21588 23278
rect 21868 23268 21924 23278
rect 21532 21698 21588 23212
rect 21756 23212 21868 23268
rect 21756 22482 21812 23212
rect 21868 23202 21924 23212
rect 21756 22430 21758 22482
rect 21810 22430 21812 22482
rect 21756 22418 21812 22430
rect 21532 21646 21534 21698
rect 21586 21646 21588 21698
rect 21532 20914 21588 21646
rect 21644 21588 21700 21626
rect 21644 21522 21700 21532
rect 21532 20862 21534 20914
rect 21586 20862 21588 20914
rect 21532 20850 21588 20862
rect 21980 20578 22036 20590
rect 21980 20526 21982 20578
rect 22034 20526 22036 20578
rect 21980 20356 22036 20526
rect 21980 20290 22036 20300
rect 21532 19124 21588 19134
rect 21420 19068 21532 19124
rect 21532 19058 21588 19068
rect 21420 18340 21476 18350
rect 21420 18246 21476 18284
rect 21532 17780 21588 17790
rect 21308 17668 21364 17678
rect 21308 17106 21364 17612
rect 21308 17054 21310 17106
rect 21362 17054 21364 17106
rect 21308 17042 21364 17054
rect 21420 16882 21476 16894
rect 21420 16830 21422 16882
rect 21474 16830 21476 16882
rect 20860 15874 21252 15876
rect 20860 15822 20862 15874
rect 20914 15822 21252 15874
rect 20860 15820 21252 15822
rect 21308 16324 21364 16334
rect 20860 15810 20916 15820
rect 20972 15316 21028 15326
rect 20972 15222 21028 15260
rect 21196 15202 21252 15214
rect 21196 15150 21198 15202
rect 21250 15150 21252 15202
rect 20748 15092 21028 15148
rect 20748 14308 20804 14318
rect 20972 14308 21028 15092
rect 21196 14868 21252 15150
rect 21196 14802 21252 14812
rect 20748 14306 20916 14308
rect 20748 14254 20750 14306
rect 20802 14254 20916 14306
rect 20748 14252 20916 14254
rect 20748 14242 20804 14252
rect 20860 14084 20916 14252
rect 20972 14242 21028 14252
rect 21196 14530 21252 14542
rect 21196 14478 21198 14530
rect 21250 14478 21252 14530
rect 21196 14084 21252 14478
rect 20860 14028 21252 14084
rect 20860 13748 20916 13758
rect 20860 13654 20916 13692
rect 20748 12180 20804 12190
rect 20636 12178 20804 12180
rect 20636 12126 20750 12178
rect 20802 12126 20804 12178
rect 20636 12124 20804 12126
rect 20748 12114 20804 12124
rect 20972 12068 21028 12078
rect 20748 11396 20804 11406
rect 20748 11302 20804 11340
rect 20972 10948 21028 12012
rect 21308 10948 21364 16268
rect 21420 15988 21476 16830
rect 21420 15922 21476 15932
rect 21420 15316 21476 15326
rect 21420 15222 21476 15260
rect 21420 14308 21476 14318
rect 21420 14214 21476 14252
rect 21532 13972 21588 17724
rect 21644 17668 21700 17678
rect 21644 16436 21700 17612
rect 21980 17444 22036 17454
rect 22092 17444 22148 26012
rect 22204 23268 22260 27580
rect 22316 27570 22372 27580
rect 22316 27300 22372 27310
rect 22540 27300 22596 35420
rect 22876 34916 22932 34954
rect 22876 34850 22932 34860
rect 22876 34692 22932 34702
rect 23100 34692 23156 40684
rect 23212 39620 23268 39630
rect 23212 38050 23268 39564
rect 23324 39618 23380 39630
rect 23324 39566 23326 39618
rect 23378 39566 23380 39618
rect 23324 38274 23380 39566
rect 23772 39508 23828 39518
rect 23772 39414 23828 39452
rect 23996 39506 24052 39518
rect 23996 39454 23998 39506
rect 24050 39454 24052 39506
rect 23660 39394 23716 39406
rect 23660 39342 23662 39394
rect 23714 39342 23716 39394
rect 23660 39060 23716 39342
rect 23660 39004 23940 39060
rect 23884 38946 23940 39004
rect 23884 38894 23886 38946
rect 23938 38894 23940 38946
rect 23884 38882 23940 38894
rect 23996 38948 24052 39454
rect 23996 38882 24052 38892
rect 24108 38668 24164 41244
rect 25228 40964 25284 40974
rect 25004 40404 25060 40414
rect 24668 38836 24724 38846
rect 24668 38668 24724 38780
rect 23324 38222 23326 38274
rect 23378 38222 23380 38274
rect 23324 38210 23380 38222
rect 23996 38612 24164 38668
rect 24556 38612 24724 38668
rect 23212 37998 23214 38050
rect 23266 37998 23268 38050
rect 23212 37986 23268 37998
rect 23212 37828 23268 37838
rect 23324 37828 23380 37838
rect 23268 37826 23380 37828
rect 23268 37774 23326 37826
rect 23378 37774 23380 37826
rect 23268 37772 23380 37774
rect 23212 34804 23268 37772
rect 23324 37762 23380 37772
rect 23548 37044 23604 37054
rect 23548 35700 23604 36988
rect 23548 35634 23604 35644
rect 23324 35588 23380 35598
rect 23324 35494 23380 35532
rect 23212 34738 23268 34748
rect 22876 34690 23156 34692
rect 22876 34638 22878 34690
rect 22930 34638 23156 34690
rect 22876 34636 23156 34638
rect 23324 34692 23380 34702
rect 22876 33460 22932 34636
rect 23100 33684 23156 33694
rect 23100 33570 23156 33628
rect 23100 33518 23102 33570
rect 23154 33518 23156 33570
rect 23100 33506 23156 33518
rect 22876 33394 22932 33404
rect 22652 33236 22708 33246
rect 22652 33122 22708 33180
rect 22988 33236 23044 33246
rect 22988 33142 23044 33180
rect 22652 33070 22654 33122
rect 22706 33070 22708 33122
rect 22652 30548 22708 33070
rect 23212 31892 23268 31902
rect 22764 31332 22820 31342
rect 22764 31218 22820 31276
rect 22764 31166 22766 31218
rect 22818 31166 22820 31218
rect 22764 31154 22820 31166
rect 23212 31220 23268 31836
rect 23212 31126 23268 31164
rect 22652 30482 22708 30492
rect 23100 27860 23156 27870
rect 22764 27858 23156 27860
rect 22764 27806 23102 27858
rect 23154 27806 23156 27858
rect 22764 27804 23156 27806
rect 22764 27746 22820 27804
rect 23100 27794 23156 27804
rect 23324 27748 23380 34636
rect 23772 34020 23828 34030
rect 23548 34018 23828 34020
rect 23548 33966 23774 34018
rect 23826 33966 23828 34018
rect 23548 33964 23828 33966
rect 23548 30548 23604 33964
rect 23772 33954 23828 33964
rect 23996 32788 24052 38612
rect 24556 35924 24612 38612
rect 24108 35922 24612 35924
rect 24108 35870 24558 35922
rect 24610 35870 24612 35922
rect 24108 35868 24612 35870
rect 24108 35698 24164 35868
rect 24108 35646 24110 35698
rect 24162 35646 24164 35698
rect 24108 35634 24164 35646
rect 24332 34914 24388 34926
rect 24332 34862 24334 34914
rect 24386 34862 24388 34914
rect 24332 33684 24388 34862
rect 24444 34356 24500 35868
rect 24556 35858 24612 35868
rect 24892 35140 24948 35150
rect 24892 35046 24948 35084
rect 24556 34914 24612 34926
rect 24556 34862 24558 34914
rect 24610 34862 24612 34914
rect 24556 34804 24612 34862
rect 24556 34738 24612 34748
rect 24444 34130 24500 34300
rect 24444 34078 24446 34130
rect 24498 34078 24500 34130
rect 24444 34066 24500 34078
rect 25004 34132 25060 40348
rect 25004 34066 25060 34076
rect 24332 33618 24388 33628
rect 25228 33460 25284 40908
rect 25340 39058 25396 41916
rect 27916 41972 27972 41982
rect 27580 41860 27636 41870
rect 25340 39006 25342 39058
rect 25394 39006 25396 39058
rect 25340 38836 25396 39006
rect 25340 38770 25396 38780
rect 26124 41188 26180 41198
rect 26124 39732 26180 41132
rect 27580 41188 27636 41804
rect 27580 41094 27636 41132
rect 27804 41074 27860 41086
rect 27804 41022 27806 41074
rect 27858 41022 27860 41074
rect 27132 40964 27188 40974
rect 26572 40740 26628 40750
rect 26572 40626 26628 40684
rect 26572 40574 26574 40626
rect 26626 40574 26628 40626
rect 26572 40562 26628 40574
rect 27020 40516 27076 40526
rect 27020 40422 27076 40460
rect 26908 40402 26964 40414
rect 26908 40350 26910 40402
rect 26962 40350 26964 40402
rect 26908 40292 26964 40350
rect 26124 39730 26628 39732
rect 26124 39678 26126 39730
rect 26178 39678 26628 39730
rect 26124 39676 26628 39678
rect 26124 38668 26180 39676
rect 26460 39506 26516 39518
rect 26460 39454 26462 39506
rect 26514 39454 26516 39506
rect 26460 39396 26516 39454
rect 26572 39506 26628 39676
rect 26908 39620 26964 40236
rect 27132 39844 27188 40908
rect 27580 40740 27636 40750
rect 27580 40514 27636 40684
rect 27804 40626 27860 41022
rect 27804 40574 27806 40626
rect 27858 40574 27860 40626
rect 27804 40562 27860 40574
rect 27580 40462 27582 40514
rect 27634 40462 27636 40514
rect 27244 40404 27300 40414
rect 27244 40402 27412 40404
rect 27244 40350 27246 40402
rect 27298 40350 27412 40402
rect 27244 40348 27412 40350
rect 27244 40338 27300 40348
rect 27132 39778 27188 39788
rect 27244 39620 27300 39630
rect 26964 39618 27300 39620
rect 26964 39566 27246 39618
rect 27298 39566 27300 39618
rect 26964 39564 27300 39566
rect 27356 39620 27412 40348
rect 27468 40402 27524 40414
rect 27468 40350 27470 40402
rect 27522 40350 27524 40402
rect 27468 39844 27524 40350
rect 27580 40404 27636 40462
rect 27580 40338 27636 40348
rect 27468 39778 27524 39788
rect 27916 39844 27972 41916
rect 28476 41972 28532 42028
rect 28476 41906 28532 41916
rect 28588 41858 28644 41870
rect 28588 41806 28590 41858
rect 28642 41806 28644 41858
rect 28588 41412 28644 41806
rect 28028 41356 28644 41412
rect 28028 41298 28084 41356
rect 28028 41246 28030 41298
rect 28082 41246 28084 41298
rect 28028 41234 28084 41246
rect 28252 41188 28308 41198
rect 28476 41188 28532 41198
rect 28252 41186 28420 41188
rect 28252 41134 28254 41186
rect 28306 41134 28420 41186
rect 28252 41132 28420 41134
rect 28252 41122 28308 41132
rect 28140 40964 28196 40974
rect 28140 40626 28196 40908
rect 28140 40574 28142 40626
rect 28194 40574 28196 40626
rect 28140 40562 28196 40574
rect 28364 40626 28420 41132
rect 28364 40574 28366 40626
rect 28418 40574 28420 40626
rect 28364 40562 28420 40574
rect 28028 40402 28084 40414
rect 28028 40350 28030 40402
rect 28082 40350 28084 40402
rect 28028 40292 28084 40350
rect 28028 40226 28084 40236
rect 27916 39778 27972 39788
rect 28140 39732 28196 39742
rect 28140 39638 28196 39676
rect 27580 39620 27636 39630
rect 27916 39620 27972 39630
rect 27356 39564 27524 39620
rect 26908 39554 26964 39564
rect 27244 39554 27300 39564
rect 26572 39454 26574 39506
rect 26626 39454 26628 39506
rect 26572 39442 26628 39454
rect 26460 39330 26516 39340
rect 26796 39394 26852 39406
rect 26796 39342 26798 39394
rect 26850 39342 26852 39394
rect 25788 38612 26180 38668
rect 26572 38724 26628 38762
rect 26572 38658 26628 38668
rect 25340 34356 25396 34366
rect 25340 34262 25396 34300
rect 25228 33394 25284 33404
rect 23996 32732 24388 32788
rect 23660 32004 23716 32014
rect 23660 31556 23716 31948
rect 23660 31490 23716 31500
rect 23436 30492 23604 30548
rect 23436 27860 23492 30492
rect 24108 30436 24164 30446
rect 23772 30100 23828 30110
rect 23660 30098 23828 30100
rect 23660 30046 23774 30098
rect 23826 30046 23828 30098
rect 23660 30044 23828 30046
rect 23436 27804 23604 27860
rect 22764 27694 22766 27746
rect 22818 27694 22820 27746
rect 22764 27634 22820 27694
rect 23212 27692 23380 27748
rect 22764 27582 22766 27634
rect 22818 27582 22820 27634
rect 22764 27570 22820 27582
rect 23100 27634 23156 27646
rect 23100 27582 23102 27634
rect 23154 27582 23156 27634
rect 22316 27206 22372 27244
rect 22428 27244 22596 27300
rect 23100 27300 23156 27582
rect 22316 27076 22372 27086
rect 22316 26982 22372 27020
rect 22428 26908 22484 27244
rect 23100 27234 23156 27244
rect 22764 27132 22932 27188
rect 22428 26852 22708 26908
rect 22540 26516 22596 26526
rect 22540 26422 22596 26460
rect 22316 25396 22372 25406
rect 22316 24946 22372 25340
rect 22316 24894 22318 24946
rect 22370 24894 22372 24946
rect 22316 24882 22372 24894
rect 22204 23202 22260 23212
rect 22428 22708 22484 22718
rect 22204 22148 22260 22158
rect 22260 22092 22372 22148
rect 22204 22082 22260 22092
rect 22204 21812 22260 21822
rect 22204 21718 22260 21756
rect 22316 21028 22372 22092
rect 22036 17388 22148 17444
rect 22204 20972 22372 21028
rect 21980 17378 22036 17388
rect 21868 16884 21924 16894
rect 21868 16790 21924 16828
rect 22204 16660 22260 20972
rect 22316 20802 22372 20814
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 22316 20356 22372 20750
rect 22316 20290 22372 20300
rect 22204 16594 22260 16604
rect 21644 16210 21700 16380
rect 21644 16158 21646 16210
rect 21698 16158 21700 16210
rect 21644 16146 21700 16158
rect 21980 15988 22036 15998
rect 21644 15428 21700 15438
rect 21644 15334 21700 15372
rect 21980 15426 22036 15932
rect 21980 15374 21982 15426
rect 22034 15374 22036 15426
rect 21980 15362 22036 15374
rect 22092 15428 22148 15438
rect 22092 14980 22148 15372
rect 22316 15316 22372 15326
rect 22316 15222 22372 15260
rect 22092 14914 22148 14924
rect 21644 14756 21700 14766
rect 21644 14530 21700 14700
rect 21644 14478 21646 14530
rect 21698 14478 21700 14530
rect 21644 14466 21700 14478
rect 21868 14532 21924 14542
rect 21868 14438 21924 14476
rect 21532 13860 21588 13916
rect 21532 13804 21700 13860
rect 21532 13636 21588 13646
rect 21532 13542 21588 13580
rect 21532 12964 21588 12974
rect 21644 12964 21700 13804
rect 21756 13746 21812 13758
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 21756 13636 21812 13694
rect 21756 13570 21812 13580
rect 21588 12908 21700 12964
rect 21756 13412 21812 13422
rect 21532 12870 21588 12908
rect 21420 12292 21476 12302
rect 21476 12236 21700 12292
rect 21420 12226 21476 12236
rect 20636 10892 21028 10948
rect 20636 10834 20692 10892
rect 20636 10782 20638 10834
rect 20690 10782 20692 10834
rect 20636 10770 20692 10782
rect 20972 10834 21028 10892
rect 20972 10782 20974 10834
rect 21026 10782 21028 10834
rect 20972 10770 21028 10782
rect 21084 10892 21364 10948
rect 21644 11618 21700 12236
rect 21644 11566 21646 11618
rect 21698 11566 21700 11618
rect 21084 10612 21140 10892
rect 21196 10724 21252 10734
rect 21644 10724 21700 11566
rect 21196 10722 21700 10724
rect 21196 10670 21198 10722
rect 21250 10670 21700 10722
rect 21196 10668 21700 10670
rect 21196 10658 21252 10668
rect 20300 9998 20302 10050
rect 20354 9998 20356 10050
rect 20300 9986 20356 9998
rect 20748 10556 21140 10612
rect 21644 10610 21700 10668
rect 21644 10558 21646 10610
rect 21698 10558 21700 10610
rect 20076 9762 20132 9772
rect 20524 9828 20580 9838
rect 20188 9716 20244 9726
rect 19628 9604 19684 9614
rect 20076 9604 20132 9642
rect 19628 9602 20076 9604
rect 19628 9550 19630 9602
rect 19682 9550 20076 9602
rect 19628 9548 20076 9550
rect 19628 9538 19684 9548
rect 20076 9538 20132 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20076 9268 20132 9278
rect 19516 9266 20132 9268
rect 19516 9214 20078 9266
rect 20130 9214 20132 9266
rect 19516 9212 20132 9214
rect 19516 9154 19572 9212
rect 20076 9202 20132 9212
rect 19516 9102 19518 9154
rect 19570 9102 19572 9154
rect 19516 9090 19572 9102
rect 20188 9156 20244 9660
rect 20188 9154 20468 9156
rect 20188 9102 20190 9154
rect 20242 9102 20468 9154
rect 20188 9100 20468 9102
rect 20188 9090 20244 9100
rect 19292 8990 19294 9042
rect 19346 8990 19348 9042
rect 19292 8978 19348 8990
rect 19740 9044 19796 9054
rect 19740 8950 19796 8988
rect 19628 8932 19684 8942
rect 19180 8866 19236 8876
rect 19516 8930 19684 8932
rect 19516 8878 19630 8930
rect 19682 8878 19684 8930
rect 19516 8876 19684 8878
rect 19516 7586 19572 8876
rect 19628 8866 19684 8876
rect 20076 8932 20132 8942
rect 20076 8370 20132 8876
rect 20076 8318 20078 8370
rect 20130 8318 20132 8370
rect 20076 8306 20132 8318
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19516 7534 19518 7586
rect 19570 7534 19572 7586
rect 19516 7522 19572 7534
rect 20412 7588 20468 9100
rect 20524 9154 20580 9772
rect 20524 9102 20526 9154
rect 20578 9102 20580 9154
rect 20524 9044 20580 9102
rect 20748 9156 20804 10556
rect 21644 10546 21700 10558
rect 20748 9062 20804 9100
rect 20860 10386 20916 10398
rect 20860 10334 20862 10386
rect 20914 10334 20916 10386
rect 20860 9044 20916 10334
rect 21756 9156 21812 13356
rect 21980 11508 22036 11518
rect 21980 11506 22372 11508
rect 21980 11454 21982 11506
rect 22034 11454 22372 11506
rect 21980 11452 22372 11454
rect 21980 11442 22036 11452
rect 21868 11396 21924 11406
rect 21868 11282 21924 11340
rect 21868 11230 21870 11282
rect 21922 11230 21924 11282
rect 21868 11218 21924 11230
rect 21868 10722 21924 10734
rect 21868 10670 21870 10722
rect 21922 10670 21924 10722
rect 21868 9828 21924 10670
rect 22316 10050 22372 11452
rect 22316 9998 22318 10050
rect 22370 9998 22372 10050
rect 22316 9986 22372 9998
rect 22428 10052 22484 22652
rect 22540 21588 22596 21598
rect 22540 21494 22596 21532
rect 22540 20804 22596 20814
rect 22540 20710 22596 20748
rect 22652 20020 22708 26852
rect 22764 26628 22820 27132
rect 22876 27074 22932 27132
rect 22876 27022 22878 27074
rect 22930 27022 22932 27074
rect 22876 27010 22932 27022
rect 22988 27020 23156 27076
rect 22988 26852 23044 27020
rect 23100 26962 23156 27020
rect 23100 26910 23102 26962
rect 23154 26910 23156 26962
rect 23100 26898 23156 26910
rect 22988 26786 23044 26796
rect 22876 26628 22932 26638
rect 22764 26572 22876 26628
rect 22876 26290 22932 26572
rect 22876 26238 22878 26290
rect 22930 26238 22932 26290
rect 22876 24836 22932 26238
rect 23100 26290 23156 26302
rect 23100 26238 23102 26290
rect 23154 26238 23156 26290
rect 23100 26068 23156 26238
rect 23100 26002 23156 26012
rect 22876 24770 22932 24780
rect 23212 25618 23268 27692
rect 23436 27636 23492 27646
rect 23436 27542 23492 27580
rect 23436 27188 23492 27198
rect 23324 27076 23380 27114
rect 23324 27010 23380 27020
rect 23436 27074 23492 27132
rect 23436 27022 23438 27074
rect 23490 27022 23492 27074
rect 23436 27010 23492 27022
rect 23548 26908 23604 27804
rect 23324 26852 23604 26908
rect 23324 26514 23380 26852
rect 23660 26850 23716 30044
rect 23772 30034 23828 30044
rect 23884 27748 23940 27758
rect 23660 26798 23662 26850
rect 23714 26798 23716 26850
rect 23660 26786 23716 26798
rect 23772 27746 23940 27748
rect 23772 27694 23886 27746
rect 23938 27694 23940 27746
rect 23772 27692 23940 27694
rect 23772 26852 23828 27692
rect 23884 27682 23940 27692
rect 23996 27636 24052 27646
rect 23996 27298 24052 27580
rect 24108 27412 24164 30380
rect 24108 27346 24164 27356
rect 23996 27246 23998 27298
rect 24050 27246 24052 27298
rect 23772 26628 23828 26796
rect 23324 26462 23326 26514
rect 23378 26462 23380 26514
rect 23324 26450 23380 26462
rect 23548 26572 23828 26628
rect 23884 27188 23940 27198
rect 23884 26964 23940 27132
rect 23436 26068 23492 26078
rect 23436 25974 23492 26012
rect 23212 25566 23214 25618
rect 23266 25566 23268 25618
rect 22652 19954 22708 19964
rect 22764 23716 22820 23726
rect 22540 16996 22596 17006
rect 22540 16902 22596 16940
rect 22652 15316 22708 15326
rect 22652 15222 22708 15260
rect 22540 14308 22596 14318
rect 22540 13858 22596 14252
rect 22540 13806 22542 13858
rect 22594 13806 22596 13858
rect 22540 13794 22596 13806
rect 21868 9734 21924 9772
rect 22204 9828 22260 9838
rect 22428 9828 22484 9996
rect 22204 9734 22260 9772
rect 22316 9826 22484 9828
rect 22316 9774 22430 9826
rect 22482 9774 22484 9826
rect 22316 9772 22484 9774
rect 22316 9380 22372 9772
rect 22428 9762 22484 9772
rect 22764 9828 22820 23660
rect 23100 22148 23156 22158
rect 22876 22092 23100 22148
rect 22876 21700 22932 22092
rect 23100 22054 23156 22092
rect 23212 21812 23268 25566
rect 23436 25732 23492 25742
rect 23324 23828 23380 23838
rect 23324 23734 23380 23772
rect 22876 21606 22932 21644
rect 23100 21756 23268 21812
rect 23324 23492 23380 23502
rect 22988 21588 23044 21598
rect 22876 21028 22932 21038
rect 22988 21028 23044 21532
rect 22876 21026 23044 21028
rect 22876 20974 22878 21026
rect 22930 20974 23044 21026
rect 22876 20972 23044 20974
rect 22876 20962 22932 20972
rect 22876 19906 22932 19918
rect 22876 19854 22878 19906
rect 22930 19854 22932 19906
rect 22876 19794 22932 19854
rect 22876 19742 22878 19794
rect 22930 19742 22932 19794
rect 22876 19684 22932 19742
rect 22876 19618 22932 19628
rect 23100 17780 23156 21756
rect 23212 21588 23268 21598
rect 23212 21494 23268 21532
rect 23324 21028 23380 23436
rect 23436 22258 23492 25676
rect 23436 22206 23438 22258
rect 23490 22206 23492 22258
rect 23436 21364 23492 22206
rect 23436 21298 23492 21308
rect 23324 20972 23492 21028
rect 23324 20804 23380 20814
rect 23212 20578 23268 20590
rect 23212 20526 23214 20578
rect 23266 20526 23268 20578
rect 23212 19794 23268 20526
rect 23212 19742 23214 19794
rect 23266 19742 23268 19794
rect 23212 19730 23268 19742
rect 23324 19906 23380 20748
rect 23436 20692 23492 20972
rect 23548 20804 23604 26572
rect 23660 26292 23716 26302
rect 23884 26292 23940 26908
rect 23660 26290 23940 26292
rect 23660 26238 23662 26290
rect 23714 26238 23940 26290
rect 23660 26236 23940 26238
rect 23660 26226 23716 26236
rect 23996 26068 24052 27246
rect 24108 27076 24164 27086
rect 24108 26982 24164 27020
rect 24332 26908 24388 32732
rect 24444 32116 24500 32126
rect 24444 31218 24500 32060
rect 24444 31166 24446 31218
rect 24498 31166 24500 31218
rect 24444 30436 24500 31166
rect 25564 31668 25620 31678
rect 24444 29988 24500 30380
rect 25228 30436 25284 30446
rect 25228 30342 25284 30380
rect 24556 30212 24612 30222
rect 24556 30118 24612 30156
rect 25004 30210 25060 30222
rect 25004 30158 25006 30210
rect 25058 30158 25060 30210
rect 24668 29988 24724 29998
rect 25004 29988 25060 30158
rect 25564 30210 25620 31612
rect 25564 30158 25566 30210
rect 25618 30158 25620 30210
rect 25564 30146 25620 30158
rect 24444 29932 24612 29988
rect 24108 26852 24164 26862
rect 24220 26852 24276 26862
rect 24332 26852 24500 26908
rect 24164 26850 24276 26852
rect 24164 26798 24222 26850
rect 24274 26798 24276 26850
rect 24164 26796 24276 26798
rect 24108 26786 24164 26796
rect 24220 26786 24276 26796
rect 24332 26516 24388 26526
rect 24332 26290 24388 26460
rect 24332 26238 24334 26290
rect 24386 26238 24388 26290
rect 23884 26066 24052 26068
rect 23884 26014 23998 26066
rect 24050 26014 24052 26066
rect 23884 26012 24052 26014
rect 23660 25844 23716 25854
rect 23660 24164 23716 25788
rect 23772 24722 23828 24734
rect 23772 24670 23774 24722
rect 23826 24670 23828 24722
rect 23772 24612 23828 24670
rect 23884 24612 23940 26012
rect 23996 26002 24052 26012
rect 24108 26178 24164 26190
rect 24108 26126 24110 26178
rect 24162 26126 24164 26178
rect 24108 26068 24164 26126
rect 24108 26002 24164 26012
rect 23996 24836 24052 24846
rect 23996 24742 24052 24780
rect 23772 24556 24276 24612
rect 23996 24276 24052 24286
rect 23884 24220 23996 24276
rect 23772 24164 23828 24174
rect 23660 24162 23828 24164
rect 23660 24110 23774 24162
rect 23826 24110 23828 24162
rect 23660 24108 23828 24110
rect 23772 24098 23828 24108
rect 23660 23826 23716 23838
rect 23660 23774 23662 23826
rect 23714 23774 23716 23826
rect 23660 22148 23716 23774
rect 23772 23828 23828 23838
rect 23772 23734 23828 23772
rect 23772 22708 23828 22718
rect 23772 22482 23828 22652
rect 23772 22430 23774 22482
rect 23826 22430 23828 22482
rect 23772 22418 23828 22430
rect 23660 22082 23716 22092
rect 23884 21810 23940 24220
rect 23996 24210 24052 24220
rect 24220 23826 24276 24556
rect 24220 23774 24222 23826
rect 24274 23774 24276 23826
rect 24220 23762 24276 23774
rect 24332 22372 24388 26238
rect 24220 22316 24388 22372
rect 24220 21924 24276 22316
rect 23884 21758 23886 21810
rect 23938 21758 23940 21810
rect 23660 21588 23716 21598
rect 23660 21494 23716 21532
rect 23884 20916 23940 21758
rect 23884 20850 23940 20860
rect 24108 21868 24276 21924
rect 24332 22146 24388 22158
rect 24332 22094 24334 22146
rect 24386 22094 24388 22146
rect 23772 20804 23828 20814
rect 23548 20802 23828 20804
rect 23548 20750 23774 20802
rect 23826 20750 23828 20802
rect 23548 20748 23828 20750
rect 23436 20636 23604 20692
rect 23324 19854 23326 19906
rect 23378 19854 23380 19906
rect 23100 17714 23156 17724
rect 23324 16436 23380 19854
rect 23324 16370 23380 16380
rect 23548 13636 23604 20636
rect 23772 20020 23828 20748
rect 23772 19954 23828 19964
rect 24108 18450 24164 21868
rect 24332 21588 24388 22094
rect 24332 21522 24388 21532
rect 24220 20916 24276 20926
rect 24220 20242 24276 20860
rect 24220 20190 24222 20242
rect 24274 20190 24276 20242
rect 24220 20178 24276 20190
rect 24444 19796 24500 26852
rect 24556 24276 24612 29932
rect 24556 24210 24612 24220
rect 24724 29932 25060 29988
rect 24668 29314 24724 29932
rect 24668 29262 24670 29314
rect 24722 29262 24724 29314
rect 24556 23826 24612 23838
rect 24556 23774 24558 23826
rect 24610 23774 24612 23826
rect 24556 22484 24612 23774
rect 24668 23828 24724 29262
rect 24780 27748 24836 27758
rect 24780 27746 25060 27748
rect 24780 27694 24782 27746
rect 24834 27694 25060 27746
rect 24780 27692 25060 27694
rect 24780 27682 24836 27692
rect 25004 27074 25060 27692
rect 25228 27746 25284 27758
rect 25228 27694 25230 27746
rect 25282 27694 25284 27746
rect 25228 27300 25284 27694
rect 25228 27244 25508 27300
rect 25004 27022 25006 27074
rect 25058 27022 25060 27074
rect 24668 23762 24724 23772
rect 24892 26964 24948 26974
rect 24892 23826 24948 26908
rect 25004 26516 25060 27022
rect 25228 27076 25284 27114
rect 25228 27010 25284 27020
rect 25340 26962 25396 26974
rect 25340 26910 25342 26962
rect 25394 26910 25396 26962
rect 25340 26908 25396 26910
rect 25004 26450 25060 26460
rect 25228 26852 25396 26908
rect 25228 25844 25284 26852
rect 25340 26786 25396 26796
rect 25452 26404 25508 27244
rect 25676 27074 25732 27086
rect 25676 27022 25678 27074
rect 25730 27022 25732 27074
rect 25676 26964 25732 27022
rect 25676 26898 25732 26908
rect 25452 26338 25508 26348
rect 25340 26178 25396 26190
rect 25340 26126 25342 26178
rect 25394 26126 25396 26178
rect 25340 25956 25396 26126
rect 25340 25890 25396 25900
rect 25228 25778 25284 25788
rect 25788 24052 25844 38612
rect 26796 38500 26852 39342
rect 26908 39396 26964 39406
rect 26908 38946 26964 39340
rect 27356 39394 27412 39406
rect 27356 39342 27358 39394
rect 27410 39342 27412 39394
rect 27356 39284 27412 39342
rect 27132 39228 27356 39284
rect 26908 38894 26910 38946
rect 26962 38894 26964 38946
rect 26908 38882 26964 38894
rect 27020 38946 27076 38958
rect 27020 38894 27022 38946
rect 27074 38894 27076 38946
rect 27020 38724 27076 38894
rect 27020 38658 27076 38668
rect 26796 38434 26852 38444
rect 27132 38052 27188 39228
rect 27356 39218 27412 39228
rect 27356 39060 27412 39070
rect 27244 39004 27356 39060
rect 27244 38946 27300 39004
rect 27356 38994 27412 39004
rect 27244 38894 27246 38946
rect 27298 38894 27300 38946
rect 27244 38882 27300 38894
rect 27468 38946 27524 39564
rect 27580 39618 27972 39620
rect 27580 39566 27582 39618
rect 27634 39566 27918 39618
rect 27970 39566 27972 39618
rect 27580 39564 27972 39566
rect 27580 39554 27636 39564
rect 27916 39554 27972 39564
rect 28252 39618 28308 39630
rect 28252 39566 28254 39618
rect 28306 39566 28308 39618
rect 27580 39172 27636 39182
rect 27580 39058 27636 39116
rect 27580 39006 27582 39058
rect 27634 39006 27636 39058
rect 27580 38994 27636 39006
rect 28252 39060 28308 39566
rect 28476 39618 28532 41132
rect 28588 40964 28644 40974
rect 28588 40870 28644 40908
rect 28476 39566 28478 39618
rect 28530 39566 28532 39618
rect 28252 38994 28308 39004
rect 28364 39060 28420 39070
rect 28476 39060 28532 39566
rect 28364 39058 28532 39060
rect 28364 39006 28366 39058
rect 28418 39006 28532 39058
rect 28364 39004 28532 39006
rect 28588 40404 28644 40414
rect 28364 38994 28420 39004
rect 28588 38948 28644 40348
rect 28812 40402 28868 40414
rect 28812 40350 28814 40402
rect 28866 40350 28868 40402
rect 28812 39844 28868 40350
rect 28812 39284 28868 39788
rect 28812 39218 28868 39228
rect 28700 39060 28756 39070
rect 28700 38966 28756 39004
rect 27468 38894 27470 38946
rect 27522 38894 27524 38946
rect 27468 38882 27524 38894
rect 28476 38892 28644 38948
rect 27692 38834 27748 38846
rect 27692 38782 27694 38834
rect 27746 38782 27748 38834
rect 27132 37986 27188 37996
rect 27356 38612 27412 38622
rect 27244 37154 27300 37166
rect 27244 37102 27246 37154
rect 27298 37102 27300 37154
rect 27244 36932 27300 37102
rect 27244 36866 27300 36876
rect 26124 34244 26180 34254
rect 26460 34244 26516 34254
rect 26180 34242 26516 34244
rect 26180 34190 26462 34242
rect 26514 34190 26516 34242
rect 26180 34188 26516 34190
rect 26124 34150 26180 34188
rect 26460 34178 26516 34188
rect 26796 34132 26852 34142
rect 26124 34020 26180 34030
rect 26012 30212 26068 30222
rect 26012 30118 26068 30156
rect 25900 27298 25956 27310
rect 25900 27246 25902 27298
rect 25954 27246 25956 27298
rect 25900 27076 25956 27246
rect 25900 27010 25956 27020
rect 25452 23996 25844 24052
rect 24892 23774 24894 23826
rect 24946 23774 24948 23826
rect 24892 23762 24948 23774
rect 25116 23938 25172 23950
rect 25116 23886 25118 23938
rect 25170 23886 25172 23938
rect 24668 23492 24724 23502
rect 24668 23378 24724 23436
rect 24668 23326 24670 23378
rect 24722 23326 24724 23378
rect 24668 23314 24724 23326
rect 24556 22428 24948 22484
rect 24668 22258 24724 22270
rect 24668 22206 24670 22258
rect 24722 22206 24724 22258
rect 24668 22148 24724 22206
rect 24668 22082 24724 22092
rect 24780 22146 24836 22158
rect 24780 22094 24782 22146
rect 24834 22094 24836 22146
rect 24668 21812 24724 21822
rect 24668 21718 24724 21756
rect 24780 21476 24836 22094
rect 24892 22148 24948 22428
rect 25004 22148 25060 22158
rect 24892 22146 25060 22148
rect 24892 22094 25006 22146
rect 25058 22094 25060 22146
rect 24892 22092 25060 22094
rect 24556 20916 24612 20926
rect 24556 20822 24612 20860
rect 24668 20132 24724 20142
rect 24780 20132 24836 21420
rect 25004 20804 25060 22092
rect 25116 21588 25172 23886
rect 25228 23492 25284 23502
rect 25228 23154 25284 23436
rect 25228 23102 25230 23154
rect 25282 23102 25284 23154
rect 25228 23090 25284 23102
rect 25228 22258 25284 22270
rect 25228 22206 25230 22258
rect 25282 22206 25284 22258
rect 25228 21924 25284 22206
rect 25228 21858 25284 21868
rect 25340 22146 25396 22158
rect 25340 22094 25342 22146
rect 25394 22094 25396 22146
rect 25340 21700 25396 22094
rect 25116 21522 25172 21532
rect 25228 21644 25340 21700
rect 25004 20738 25060 20748
rect 25004 20580 25060 20590
rect 25228 20580 25284 21644
rect 25340 21634 25396 21644
rect 25340 21476 25396 21486
rect 25340 21382 25396 21420
rect 25340 20802 25396 20814
rect 25340 20750 25342 20802
rect 25394 20750 25396 20802
rect 25340 20580 25396 20750
rect 25060 20524 25396 20580
rect 25004 20486 25060 20524
rect 25452 20356 25508 23996
rect 25564 23828 25620 23838
rect 25564 23266 25620 23772
rect 25564 23214 25566 23266
rect 25618 23214 25620 23266
rect 25564 23202 25620 23214
rect 25788 23042 25844 23054
rect 25788 22990 25790 23042
rect 25842 22990 25844 23042
rect 25564 22148 25620 22158
rect 25564 22054 25620 22092
rect 24724 20076 24836 20132
rect 25340 20300 25508 20356
rect 25564 20916 25620 20926
rect 24668 20038 24724 20076
rect 24556 19796 24612 19806
rect 24444 19740 24556 19796
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 23548 13570 23604 13580
rect 23772 18340 23828 18350
rect 24108 18340 24164 18398
rect 23772 18338 24164 18340
rect 23772 18286 23774 18338
rect 23826 18286 24164 18338
rect 23772 18284 24164 18286
rect 24556 18338 24612 19740
rect 25340 18452 25396 20300
rect 25452 20132 25508 20142
rect 25452 20018 25508 20076
rect 25452 19966 25454 20018
rect 25506 19966 25508 20018
rect 25452 19954 25508 19966
rect 25564 20020 25620 20860
rect 25676 20020 25732 20030
rect 25564 20018 25732 20020
rect 25564 19966 25678 20018
rect 25730 19966 25732 20018
rect 25564 19964 25732 19966
rect 25676 19954 25732 19964
rect 25676 19124 25732 19134
rect 25676 18674 25732 19068
rect 25676 18622 25678 18674
rect 25730 18622 25732 18674
rect 25676 18610 25732 18622
rect 25340 18396 25732 18452
rect 24556 18286 24558 18338
rect 24610 18286 24612 18338
rect 23548 12962 23604 12974
rect 23548 12910 23550 12962
rect 23602 12910 23604 12962
rect 23548 11844 23604 12910
rect 23548 11778 23604 11788
rect 23660 12740 23716 12750
rect 23660 11508 23716 12684
rect 23772 12068 23828 18284
rect 24556 18004 24612 18286
rect 24556 17938 24612 17948
rect 25340 18116 25396 18126
rect 25340 17778 25396 18060
rect 25340 17726 25342 17778
rect 25394 17726 25396 17778
rect 25340 17714 25396 17726
rect 25676 17778 25732 18396
rect 25676 17726 25678 17778
rect 25730 17726 25732 17778
rect 25676 17668 25732 17726
rect 25676 17602 25732 17612
rect 25004 17220 25060 17230
rect 24668 17108 24724 17118
rect 24668 16770 24724 17052
rect 24668 16718 24670 16770
rect 24722 16718 24724 16770
rect 24668 16706 24724 16718
rect 24220 14868 24276 14878
rect 24220 13074 24276 14812
rect 24668 13636 24724 13646
rect 24668 13542 24724 13580
rect 24220 13022 24222 13074
rect 24274 13022 24276 13074
rect 24220 13010 24276 13022
rect 23772 12002 23828 12012
rect 23660 11442 23716 11452
rect 25004 10164 25060 17164
rect 25452 16884 25508 16894
rect 25228 16548 25284 16558
rect 25228 15652 25284 16492
rect 25228 15586 25284 15596
rect 25452 11844 25508 16828
rect 25788 15148 25844 22990
rect 25900 22146 25956 22158
rect 25900 22094 25902 22146
rect 25954 22094 25956 22146
rect 25900 21700 25956 22094
rect 26124 21924 26180 33964
rect 26236 33460 26292 33470
rect 26236 28420 26292 33404
rect 26572 32788 26628 32798
rect 26796 32788 26852 34076
rect 26908 34132 26964 34142
rect 26908 34018 26964 34076
rect 26908 33966 26910 34018
rect 26962 33966 26964 34018
rect 26908 33954 26964 33966
rect 27356 33796 27412 38556
rect 27692 38500 27748 38782
rect 27916 38836 27972 38874
rect 27916 38770 27972 38780
rect 28252 38724 28308 38734
rect 28476 38668 28532 38892
rect 27692 38434 27748 38444
rect 27916 38612 27972 38622
rect 27916 37492 27972 38556
rect 27916 37378 27972 37436
rect 27916 37326 27918 37378
rect 27970 37326 27972 37378
rect 27916 37314 27972 37326
rect 28140 37378 28196 37390
rect 28140 37326 28142 37378
rect 28194 37326 28196 37378
rect 28140 36932 28196 37326
rect 27468 34020 27524 34030
rect 27468 34018 27636 34020
rect 27468 33966 27470 34018
rect 27522 33966 27636 34018
rect 27468 33964 27636 33966
rect 27468 33954 27524 33964
rect 26908 33740 27412 33796
rect 26908 32900 26964 33740
rect 27020 33460 27076 33470
rect 27580 33460 27636 33964
rect 27076 33404 27524 33460
rect 27020 33366 27076 33404
rect 26908 32834 26964 32844
rect 27356 33234 27412 33246
rect 27356 33182 27358 33234
rect 27410 33182 27412 33234
rect 26572 32786 26796 32788
rect 26572 32734 26574 32786
rect 26626 32734 26796 32786
rect 26572 32732 26796 32734
rect 26572 32722 26628 32732
rect 26796 32722 26852 32732
rect 26908 32676 26964 32686
rect 27020 32676 27076 32686
rect 26964 32674 27076 32676
rect 26964 32622 27022 32674
rect 27074 32622 27076 32674
rect 26964 32620 27076 32622
rect 26908 32116 26964 32620
rect 27020 32610 27076 32620
rect 27132 32564 27188 32574
rect 27356 32564 27412 33182
rect 27468 33234 27524 33404
rect 27580 33394 27636 33404
rect 28028 33460 28084 33470
rect 27692 33348 27748 33358
rect 27692 33254 27748 33292
rect 27916 33236 27972 33246
rect 27468 33182 27470 33234
rect 27522 33182 27524 33234
rect 27468 33170 27524 33182
rect 27804 33234 27972 33236
rect 27804 33182 27918 33234
rect 27970 33182 27972 33234
rect 27804 33180 27972 33182
rect 27804 32900 27860 33180
rect 27916 33170 27972 33180
rect 28028 33234 28084 33404
rect 28028 33182 28030 33234
rect 28082 33182 28084 33234
rect 28028 33170 28084 33182
rect 27132 32562 27412 32564
rect 27132 32510 27134 32562
rect 27186 32510 27412 32562
rect 27132 32508 27412 32510
rect 27468 32844 27860 32900
rect 27468 32674 27524 32844
rect 27468 32622 27470 32674
rect 27522 32622 27524 32674
rect 27020 32452 27076 32462
rect 27020 32338 27076 32396
rect 27020 32286 27022 32338
rect 27074 32286 27076 32338
rect 27020 32274 27076 32286
rect 26908 32060 27076 32116
rect 26908 31444 26964 31454
rect 26684 29316 26740 29326
rect 26236 28354 26292 28364
rect 26460 28644 26516 28654
rect 26684 28644 26740 29260
rect 26908 28868 26964 31388
rect 26236 27300 26292 27310
rect 26236 27074 26292 27244
rect 26348 27188 26404 27198
rect 26348 27094 26404 27132
rect 26236 27022 26238 27074
rect 26290 27022 26292 27074
rect 26236 27010 26292 27022
rect 26460 27074 26516 28588
rect 26460 27022 26462 27074
rect 26514 27022 26516 27074
rect 26460 27010 26516 27022
rect 26572 28642 26740 28644
rect 26572 28590 26686 28642
rect 26738 28590 26740 28642
rect 26572 28588 26740 28590
rect 26572 26852 26628 28588
rect 26684 28578 26740 28588
rect 26796 28812 26964 28868
rect 26572 26786 26628 26796
rect 26684 28420 26740 28430
rect 26124 21858 26180 21868
rect 26348 24836 26404 24846
rect 25900 21634 25956 21644
rect 26236 20804 26292 20814
rect 25900 20578 25956 20590
rect 25900 20526 25902 20578
rect 25954 20526 25956 20578
rect 25900 19908 25956 20526
rect 25900 19842 25956 19852
rect 26012 19794 26068 19806
rect 26012 19742 26014 19794
rect 26066 19742 26068 19794
rect 26012 17444 26068 19742
rect 26124 18116 26180 18126
rect 26124 17666 26180 18060
rect 26124 17614 26126 17666
rect 26178 17614 26180 17666
rect 26124 17602 26180 17614
rect 26012 17378 26068 17388
rect 26012 15652 26068 15662
rect 26012 15538 26068 15596
rect 26012 15486 26014 15538
rect 26066 15486 26068 15538
rect 26012 15474 26068 15486
rect 26236 15148 26292 20748
rect 26348 20130 26404 24780
rect 26684 20244 26740 28364
rect 26796 27300 26852 28812
rect 26908 28644 26964 28654
rect 26908 28530 26964 28588
rect 26908 28478 26910 28530
rect 26962 28478 26964 28530
rect 26908 28466 26964 28478
rect 26908 27300 26964 27310
rect 26796 27244 26908 27300
rect 26908 27206 26964 27244
rect 26796 26962 26852 26974
rect 26796 26910 26798 26962
rect 26850 26910 26852 26962
rect 26796 26404 26852 26910
rect 27020 26908 27076 32060
rect 27132 31668 27188 32508
rect 27244 31668 27300 31678
rect 27132 31612 27244 31668
rect 27244 31574 27300 31612
rect 27468 31332 27524 32622
rect 27580 32674 27636 32686
rect 27580 32622 27582 32674
rect 27634 32622 27636 32674
rect 27580 31780 27636 32622
rect 27804 32564 27860 32574
rect 28028 32564 28084 32574
rect 27804 32562 28084 32564
rect 27804 32510 27806 32562
rect 27858 32510 28030 32562
rect 28082 32510 28084 32562
rect 27804 32508 28084 32510
rect 27804 32498 27860 32508
rect 28028 32498 28084 32508
rect 28140 32340 28196 36876
rect 28252 34020 28308 38668
rect 28252 33954 28308 33964
rect 28364 38612 28532 38668
rect 28364 33684 28420 38612
rect 28812 37492 28868 37502
rect 28924 37492 28980 42924
rect 29036 42532 29092 43372
rect 29260 43314 29316 43326
rect 29260 43262 29262 43314
rect 29314 43262 29316 43314
rect 29260 42756 29316 43262
rect 29372 42980 29428 44270
rect 29932 44322 29988 44334
rect 29932 44270 29934 44322
rect 29986 44270 29988 44322
rect 29932 43762 29988 44270
rect 29932 43710 29934 43762
rect 29986 43710 29988 43762
rect 29932 43698 29988 43710
rect 29596 43540 29652 43550
rect 29596 43446 29652 43484
rect 29932 43428 29988 43438
rect 30044 43428 30100 44940
rect 30156 44930 30212 44940
rect 30828 44548 30884 44558
rect 30828 44454 30884 44492
rect 30604 44212 30660 44222
rect 29988 43372 30100 43428
rect 30156 43538 30212 43550
rect 30156 43486 30158 43538
rect 30210 43486 30212 43538
rect 29932 43362 29988 43372
rect 29372 42914 29428 42924
rect 29260 42690 29316 42700
rect 29036 42196 29092 42476
rect 29260 42532 29316 42542
rect 29260 42438 29316 42476
rect 29036 42140 29316 42196
rect 29148 40628 29204 40638
rect 29148 40068 29204 40572
rect 29148 40002 29204 40012
rect 28812 37490 28980 37492
rect 28812 37438 28814 37490
rect 28866 37438 28980 37490
rect 28812 37436 28980 37438
rect 29148 38500 29204 38510
rect 29148 37826 29204 38444
rect 29148 37774 29150 37826
rect 29202 37774 29204 37826
rect 28812 37426 28868 37436
rect 28476 37268 28532 37278
rect 28476 37174 28532 37212
rect 28588 36258 28644 36270
rect 28588 36206 28590 36258
rect 28642 36206 28644 36258
rect 28588 35140 28644 36206
rect 29148 35364 29204 37774
rect 28588 35074 28644 35084
rect 28700 35308 29204 35364
rect 28588 34468 28644 34478
rect 28476 33684 28532 33694
rect 28364 33628 28476 33684
rect 28476 33618 28532 33628
rect 28588 33460 28644 34412
rect 28588 33366 28644 33404
rect 28252 33236 28308 33246
rect 28252 33142 28308 33180
rect 28364 32788 28420 32798
rect 28364 32786 28532 32788
rect 28364 32734 28366 32786
rect 28418 32734 28532 32786
rect 28364 32732 28532 32734
rect 28364 32722 28420 32732
rect 28364 32562 28420 32574
rect 28364 32510 28366 32562
rect 28418 32510 28420 32562
rect 28364 32452 28420 32510
rect 28364 32386 28420 32396
rect 27916 32284 28196 32340
rect 27580 31714 27636 31724
rect 27804 32004 27860 32014
rect 27580 31556 27636 31566
rect 27580 31462 27636 31500
rect 27244 31276 27524 31332
rect 27244 31106 27300 31276
rect 27244 31054 27246 31106
rect 27298 31054 27300 31106
rect 27244 28644 27300 31054
rect 27356 31108 27412 31118
rect 27356 31014 27412 31052
rect 27580 31108 27636 31118
rect 27580 31106 27748 31108
rect 27580 31054 27582 31106
rect 27634 31054 27748 31106
rect 27580 31052 27748 31054
rect 27580 31042 27636 31052
rect 27692 30994 27748 31052
rect 27692 30942 27694 30994
rect 27746 30942 27748 30994
rect 27692 30930 27748 30942
rect 27692 30212 27748 30222
rect 27692 29652 27748 30156
rect 27692 29426 27748 29596
rect 27692 29374 27694 29426
rect 27746 29374 27748 29426
rect 27692 29362 27748 29374
rect 27244 28578 27300 28588
rect 27580 27860 27636 27870
rect 27356 27748 27412 27758
rect 27356 27746 27524 27748
rect 27356 27694 27358 27746
rect 27410 27694 27524 27746
rect 27356 27692 27524 27694
rect 27356 27682 27412 27692
rect 27356 27300 27412 27310
rect 27356 27186 27412 27244
rect 27356 27134 27358 27186
rect 27410 27134 27412 27186
rect 27356 27122 27412 27134
rect 27468 27188 27524 27692
rect 27468 27122 27524 27132
rect 26796 26338 26852 26348
rect 26908 26852 27076 26908
rect 26796 25506 26852 25518
rect 26796 25454 26798 25506
rect 26850 25454 26852 25506
rect 26796 25284 26852 25454
rect 26796 25218 26852 25228
rect 26572 20188 26740 20244
rect 26796 24836 26852 24846
rect 26348 20078 26350 20130
rect 26402 20078 26404 20130
rect 26348 20066 26404 20078
rect 26460 20132 26516 20142
rect 26460 19124 26516 20076
rect 26460 19058 26516 19068
rect 25788 15092 26068 15148
rect 25452 11778 25508 11788
rect 25676 14308 25732 14318
rect 25676 11396 25732 14252
rect 25676 11330 25732 11340
rect 25004 10098 25060 10108
rect 23100 10052 23156 10062
rect 23100 9938 23156 9996
rect 23100 9886 23102 9938
rect 23154 9886 23156 9938
rect 23100 9874 23156 9886
rect 22764 9762 22820 9772
rect 23548 9828 23604 9838
rect 23548 9734 23604 9772
rect 24332 9828 24388 9838
rect 24332 9734 24388 9772
rect 24444 9716 24500 9726
rect 24444 9622 24500 9660
rect 25900 9716 25956 9726
rect 21644 9100 21812 9156
rect 21868 9324 22372 9380
rect 22652 9602 22708 9614
rect 22652 9550 22654 9602
rect 22706 9550 22708 9602
rect 20972 9044 21028 9054
rect 20860 9042 21028 9044
rect 20860 8990 20974 9042
rect 21026 8990 21028 9042
rect 20860 8988 21028 8990
rect 20524 8978 20580 8988
rect 20972 8978 21028 8988
rect 21308 9044 21364 9054
rect 21308 8950 21364 8988
rect 20636 8930 20692 8942
rect 20636 8878 20638 8930
rect 20690 8878 20692 8930
rect 20636 7700 20692 8878
rect 21084 7700 21140 7710
rect 20636 7644 20916 7700
rect 20412 7532 20692 7588
rect 20188 7474 20244 7486
rect 20188 7422 20190 7474
rect 20242 7422 20244 7474
rect 20188 6692 20244 7422
rect 20412 6802 20468 7532
rect 20636 7474 20692 7532
rect 20636 7422 20638 7474
rect 20690 7422 20692 7474
rect 20636 7410 20692 7422
rect 20412 6750 20414 6802
rect 20466 6750 20468 6802
rect 20412 6738 20468 6750
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19740 6132 19796 6142
rect 20188 6132 20244 6636
rect 19740 6130 20244 6132
rect 19740 6078 19742 6130
rect 19794 6078 20244 6130
rect 19740 6076 20244 6078
rect 19740 6066 19796 6076
rect 20188 5906 20244 6076
rect 20860 6018 20916 7644
rect 21084 7474 21140 7644
rect 21084 7422 21086 7474
rect 21138 7422 21140 7474
rect 21084 7410 21140 7422
rect 20860 5966 20862 6018
rect 20914 5966 20916 6018
rect 20860 5954 20916 5966
rect 21308 7250 21364 7262
rect 21308 7198 21310 7250
rect 21362 7198 21364 7250
rect 20188 5854 20190 5906
rect 20242 5854 20244 5906
rect 20188 5842 20244 5854
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19292 4114 19348 4126
rect 19292 4062 19294 4114
rect 19346 4062 19348 4114
rect 17836 3490 17892 3500
rect 19180 3556 19236 3594
rect 19180 3490 19236 3500
rect 19292 3388 19348 4062
rect 20860 3668 20916 3678
rect 20076 3556 20132 3566
rect 20076 3462 20132 3500
rect 16940 3332 17332 3388
rect 18844 3332 19348 3388
rect 16940 980 16996 3332
rect 16828 924 16996 980
rect 16828 800 16884 924
rect 18844 800 18900 3332
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 3612
rect 21308 3554 21364 7198
rect 21644 4564 21700 9100
rect 21868 9044 21924 9324
rect 22204 9156 22260 9166
rect 22260 9100 22484 9156
rect 22204 9062 22260 9100
rect 21756 8932 21812 8942
rect 21868 8932 21924 8988
rect 21756 8930 21924 8932
rect 21756 8878 21758 8930
rect 21810 8878 21924 8930
rect 21756 8876 21924 8878
rect 21756 8866 21812 8876
rect 21868 7700 21924 7710
rect 21868 7606 21924 7644
rect 22428 6916 22484 9100
rect 22652 8372 22708 9550
rect 25900 9044 25956 9660
rect 25788 9042 25956 9044
rect 25788 8990 25902 9042
rect 25954 8990 25956 9042
rect 25788 8988 25956 8990
rect 22652 8306 22708 8316
rect 23660 8372 23716 8382
rect 23660 8278 23716 8316
rect 25788 8370 25844 8988
rect 25900 8978 25956 8988
rect 25788 8318 25790 8370
rect 25842 8318 25844 8370
rect 25788 8306 25844 8318
rect 22988 8260 23044 8270
rect 22988 8166 23044 8204
rect 22652 6916 22708 6926
rect 23436 6916 23492 6926
rect 22428 6914 23492 6916
rect 22428 6862 22654 6914
rect 22706 6862 23438 6914
rect 23490 6862 23492 6914
rect 22428 6860 23492 6862
rect 22428 6802 22484 6860
rect 22652 6850 22708 6860
rect 23436 6850 23492 6860
rect 22428 6750 22430 6802
rect 22482 6750 22484 6802
rect 22428 6738 22484 6750
rect 23660 6692 23716 6702
rect 23660 6598 23716 6636
rect 24220 6692 24276 6702
rect 24220 6598 24276 6636
rect 22764 6580 22820 6590
rect 22764 6578 23044 6580
rect 22764 6526 22766 6578
rect 22818 6526 23044 6578
rect 22764 6524 23044 6526
rect 22764 6514 22820 6524
rect 22988 5794 23044 6524
rect 22988 5742 22990 5794
rect 23042 5742 23044 5794
rect 22988 5730 23044 5742
rect 23100 6466 23156 6478
rect 23100 6414 23102 6466
rect 23154 6414 23156 6466
rect 23100 5572 23156 6414
rect 22540 5516 23156 5572
rect 22540 5122 22596 5516
rect 22540 5070 22542 5122
rect 22594 5070 22596 5122
rect 22540 5058 22596 5070
rect 22652 5236 22708 5246
rect 22092 4564 22148 4574
rect 21644 4562 22148 4564
rect 21644 4510 22094 4562
rect 22146 4510 22148 4562
rect 21644 4508 22148 4510
rect 21644 4338 21700 4508
rect 22092 4498 22148 4508
rect 21644 4286 21646 4338
rect 21698 4286 21700 4338
rect 21644 4274 21700 4286
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 21308 3502 21310 3554
rect 21362 3502 21364 3554
rect 21308 3490 21364 3502
rect 22652 2436 22708 5180
rect 24108 5236 24164 5246
rect 24108 5142 24164 5180
rect 23100 5124 23156 5134
rect 22764 5122 23156 5124
rect 22764 5070 23102 5122
rect 23154 5070 23156 5122
rect 22764 5068 23156 5070
rect 22764 5010 22820 5068
rect 23100 5058 23156 5068
rect 22764 4958 22766 5010
rect 22818 4958 22820 5010
rect 22764 4946 22820 4958
rect 25340 3666 25396 3678
rect 25340 3614 25342 3666
rect 25394 3614 25396 3666
rect 25340 3388 25396 3614
rect 26012 3556 26068 15092
rect 26124 15092 26292 15148
rect 26460 15204 26516 15242
rect 26572 15204 26628 20188
rect 26684 20018 26740 20030
rect 26684 19966 26686 20018
rect 26738 19966 26740 20018
rect 26684 19236 26740 19966
rect 26796 20020 26852 24780
rect 26796 19954 26852 19964
rect 26796 19236 26852 19246
rect 26684 19234 26852 19236
rect 26684 19182 26798 19234
rect 26850 19182 26852 19234
rect 26684 19180 26852 19182
rect 26796 19170 26852 19180
rect 26908 17892 26964 26852
rect 27244 25284 27300 25294
rect 27244 25190 27300 25228
rect 27580 24610 27636 27804
rect 27580 24558 27582 24610
rect 27634 24558 27636 24610
rect 27580 24546 27636 24558
rect 27580 23940 27636 23950
rect 27580 23378 27636 23884
rect 27580 23326 27582 23378
rect 27634 23326 27636 23378
rect 27580 23314 27636 23326
rect 27692 23266 27748 23278
rect 27692 23214 27694 23266
rect 27746 23214 27748 23266
rect 27132 23156 27188 23166
rect 27692 23156 27748 23214
rect 27132 23154 27692 23156
rect 27132 23102 27134 23154
rect 27186 23102 27692 23154
rect 27132 23100 27692 23102
rect 27132 23090 27188 23100
rect 27692 23062 27748 23100
rect 27468 22930 27524 22942
rect 27468 22878 27470 22930
rect 27522 22878 27524 22930
rect 27468 22148 27524 22878
rect 27468 22082 27524 22092
rect 27020 20132 27076 20142
rect 27020 20038 27076 20076
rect 27804 19460 27860 31948
rect 27916 30996 27972 32284
rect 28364 32228 28420 32238
rect 28028 31220 28084 31230
rect 28028 31218 28308 31220
rect 28028 31166 28030 31218
rect 28082 31166 28308 31218
rect 28028 31164 28308 31166
rect 28028 31154 28084 31164
rect 28140 30996 28196 31006
rect 27916 30940 28084 30996
rect 27020 19404 27860 19460
rect 27916 28644 27972 28654
rect 27020 18788 27076 19404
rect 27916 19346 27972 28588
rect 28028 26908 28084 30940
rect 28140 30902 28196 30940
rect 28252 29540 28308 31164
rect 28364 31106 28420 32172
rect 28364 31054 28366 31106
rect 28418 31054 28420 31106
rect 28364 31042 28420 31054
rect 28476 30324 28532 32732
rect 28700 32562 28756 35308
rect 29260 35028 29316 42140
rect 30156 41188 30212 43486
rect 30492 41412 30548 41422
rect 30156 41132 30436 41188
rect 30156 39732 30212 39742
rect 30156 39638 30212 39676
rect 29484 39620 29540 39630
rect 29484 39526 29540 39564
rect 29372 39060 29428 39070
rect 29372 38052 29428 39004
rect 30380 39058 30436 41132
rect 30380 39006 30382 39058
rect 30434 39006 30436 39058
rect 30380 38994 30436 39006
rect 29372 38050 30212 38052
rect 29372 37998 29374 38050
rect 29426 37998 30212 38050
rect 29372 37996 30212 37998
rect 29372 37986 29428 37996
rect 29372 37492 29428 37502
rect 29372 37398 29428 37436
rect 29932 37268 29988 37278
rect 29932 37174 29988 37212
rect 30044 36482 30100 36494
rect 30044 36430 30046 36482
rect 30098 36430 30100 36482
rect 28700 32510 28702 32562
rect 28754 32510 28756 32562
rect 28700 32228 28756 32510
rect 28700 32162 28756 32172
rect 28812 34972 29316 35028
rect 29820 35586 29876 35598
rect 29820 35534 29822 35586
rect 29874 35534 29876 35586
rect 29820 35028 29876 35534
rect 30044 35140 30100 36430
rect 30044 35074 30100 35084
rect 28812 31892 28868 34972
rect 29148 34804 29204 34814
rect 29148 34710 29204 34748
rect 29708 34804 29764 34814
rect 29708 34710 29764 34748
rect 29260 34690 29316 34702
rect 29260 34638 29262 34690
rect 29314 34638 29316 34690
rect 29260 34244 29316 34638
rect 29820 34468 29876 34972
rect 29820 34402 29876 34412
rect 30044 34914 30100 34926
rect 30044 34862 30046 34914
rect 30098 34862 30100 34914
rect 30044 34244 30100 34862
rect 29260 34188 30100 34244
rect 29596 34020 29652 34030
rect 29260 34018 29652 34020
rect 29260 33966 29598 34018
rect 29650 33966 29652 34018
rect 29260 33964 29652 33966
rect 29148 33572 29204 33582
rect 29036 33346 29092 33358
rect 29036 33294 29038 33346
rect 29090 33294 29092 33346
rect 29036 33236 29092 33294
rect 29036 33170 29092 33180
rect 29148 32674 29204 33516
rect 29260 33458 29316 33964
rect 29596 33954 29652 33964
rect 29260 33406 29262 33458
rect 29314 33406 29316 33458
rect 29260 33394 29316 33406
rect 29484 33796 29540 33806
rect 29708 33796 29764 34188
rect 29372 33348 29428 33358
rect 29372 33254 29428 33292
rect 29372 32788 29428 32798
rect 29484 32788 29540 33740
rect 29372 32786 29540 32788
rect 29372 32734 29374 32786
rect 29426 32734 29540 32786
rect 29372 32732 29540 32734
rect 29596 33740 29764 33796
rect 29372 32722 29428 32732
rect 29148 32622 29150 32674
rect 29202 32622 29204 32674
rect 28700 31836 28868 31892
rect 29036 32562 29092 32574
rect 29036 32510 29038 32562
rect 29090 32510 29092 32562
rect 28588 30996 28644 31006
rect 28588 30902 28644 30940
rect 28476 30258 28532 30268
rect 28476 29652 28532 29662
rect 28364 29540 28420 29550
rect 28252 29538 28420 29540
rect 28252 29486 28366 29538
rect 28418 29486 28420 29538
rect 28252 29484 28420 29486
rect 28364 29474 28420 29484
rect 28476 28084 28532 29596
rect 28588 28084 28644 28094
rect 28140 28082 28644 28084
rect 28140 28030 28590 28082
rect 28642 28030 28644 28082
rect 28140 28028 28644 28030
rect 28140 27858 28196 28028
rect 28588 28018 28644 28028
rect 28140 27806 28142 27858
rect 28194 27806 28196 27858
rect 28140 27794 28196 27806
rect 28028 26852 28532 26908
rect 27916 19294 27918 19346
rect 27970 19294 27972 19346
rect 27916 19236 27972 19294
rect 27468 19180 27972 19236
rect 28028 23156 28084 23166
rect 27244 19122 27300 19134
rect 27468 19124 27524 19180
rect 27244 19070 27246 19122
rect 27298 19070 27300 19122
rect 27132 19012 27188 19022
rect 27132 18918 27188 18956
rect 27020 18732 27188 18788
rect 26908 17780 26964 17836
rect 27020 17780 27076 17790
rect 26908 17778 27076 17780
rect 26908 17726 27022 17778
rect 27074 17726 27076 17778
rect 26908 17724 27076 17726
rect 27020 17714 27076 17724
rect 26796 15652 26852 15662
rect 26796 15314 26852 15596
rect 26796 15262 26798 15314
rect 26850 15262 26852 15314
rect 26796 15250 26852 15262
rect 26516 15148 26628 15204
rect 26460 15138 26516 15148
rect 26124 14530 26180 15092
rect 27132 14644 27188 18732
rect 27244 17666 27300 19070
rect 27244 17614 27246 17666
rect 27298 17614 27300 17666
rect 27244 17602 27300 17614
rect 27356 19122 27524 19124
rect 27356 19070 27470 19122
rect 27522 19070 27524 19122
rect 27356 19068 27524 19070
rect 27132 14550 27188 14588
rect 26124 14478 26126 14530
rect 26178 14478 26180 14530
rect 26124 14466 26180 14478
rect 26348 14306 26404 14318
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 26348 13524 26404 14254
rect 26684 14308 26740 14318
rect 26684 14214 26740 14252
rect 26348 13458 26404 13468
rect 26460 14196 26516 14206
rect 26348 13076 26404 13086
rect 26460 13076 26516 14140
rect 27244 14196 27300 14206
rect 27244 13970 27300 14140
rect 27244 13918 27246 13970
rect 27298 13918 27300 13970
rect 27244 13906 27300 13918
rect 26348 13074 26516 13076
rect 26348 13022 26350 13074
rect 26402 13022 26516 13074
rect 26348 13020 26516 13022
rect 26348 13010 26404 13020
rect 27244 12852 27300 12862
rect 26796 12738 26852 12750
rect 26796 12686 26798 12738
rect 26850 12686 26852 12738
rect 26348 11844 26404 11854
rect 26236 10836 26292 10846
rect 26236 10742 26292 10780
rect 26236 9042 26292 9054
rect 26236 8990 26238 9042
rect 26290 8990 26292 9042
rect 26236 8932 26292 8990
rect 26236 8866 26292 8876
rect 26348 8260 26404 11788
rect 26796 11844 26852 12686
rect 26796 11778 26852 11788
rect 26908 11172 26964 11182
rect 26908 10052 26964 11116
rect 27244 10836 27300 12796
rect 27356 12180 27412 19068
rect 27468 19058 27524 19068
rect 27580 19012 27636 19022
rect 27636 18956 27972 19012
rect 27580 18946 27636 18956
rect 27916 18562 27972 18956
rect 27916 18510 27918 18562
rect 27970 18510 27972 18562
rect 27916 18498 27972 18510
rect 27468 17892 27524 17902
rect 27468 17554 27524 17836
rect 27468 17502 27470 17554
rect 27522 17502 27524 17554
rect 27468 17490 27524 17502
rect 27580 17556 27636 17566
rect 27580 17462 27636 17500
rect 28028 17332 28084 23100
rect 28252 23156 28308 23166
rect 28252 23062 28308 23100
rect 27804 17276 28084 17332
rect 28140 17556 28196 17566
rect 28196 17500 28308 17556
rect 27804 15652 27860 17276
rect 28140 16100 28196 17500
rect 28252 17442 28308 17500
rect 28252 17390 28254 17442
rect 28306 17390 28308 17442
rect 28252 17378 28308 17390
rect 27580 14530 27636 14542
rect 27580 14478 27582 14530
rect 27634 14478 27636 14530
rect 27580 14196 27636 14478
rect 27580 14130 27636 14140
rect 27804 13972 27860 15596
rect 27916 16044 28196 16100
rect 27916 15204 27972 16044
rect 27916 14308 27972 15148
rect 28028 15316 28084 15326
rect 28028 14530 28084 15260
rect 28476 15148 28532 26852
rect 28588 24052 28644 24062
rect 28588 23958 28644 23996
rect 28700 23042 28756 31836
rect 29036 31668 29092 32510
rect 29148 32116 29204 32622
rect 29148 32050 29204 32060
rect 29484 32338 29540 32350
rect 29484 32286 29486 32338
rect 29538 32286 29540 32338
rect 28700 22990 28702 23042
rect 28754 22990 28756 23042
rect 28588 20580 28644 20590
rect 28700 20580 28756 22990
rect 28812 31106 28868 31118
rect 28812 31054 28814 31106
rect 28866 31054 28868 31106
rect 28812 30772 28868 31054
rect 28924 31108 28980 31118
rect 29036 31108 29092 31612
rect 28924 31106 29092 31108
rect 28924 31054 28926 31106
rect 28978 31054 29092 31106
rect 28924 31052 29092 31054
rect 28924 31042 28980 31052
rect 29372 30882 29428 30894
rect 29372 30830 29374 30882
rect 29426 30830 29428 30882
rect 29372 30772 29428 30830
rect 28812 30716 29428 30772
rect 28812 23044 28868 30716
rect 29484 28644 29540 32286
rect 29148 28642 29540 28644
rect 29148 28590 29486 28642
rect 29538 28590 29540 28642
rect 29148 28588 29540 28590
rect 29148 28082 29204 28588
rect 29484 28578 29540 28588
rect 29148 28030 29150 28082
rect 29202 28030 29204 28082
rect 29148 28018 29204 28030
rect 29372 27858 29428 27870
rect 29372 27806 29374 27858
rect 29426 27806 29428 27858
rect 29372 27748 29428 27806
rect 29372 27682 29428 27692
rect 29484 26292 29540 26302
rect 29484 25618 29540 26236
rect 29484 25566 29486 25618
rect 29538 25566 29540 25618
rect 29484 25554 29540 25566
rect 29148 24052 29204 24062
rect 29148 23938 29204 23996
rect 29148 23886 29150 23938
rect 29202 23886 29204 23938
rect 29148 23874 29204 23886
rect 29484 23940 29540 23950
rect 29484 23846 29540 23884
rect 29596 23938 29652 33740
rect 30156 33348 30212 37996
rect 30492 35252 30548 41356
rect 30492 35186 30548 35196
rect 30604 35138 30660 44156
rect 31612 43652 31668 43662
rect 31612 43558 31668 43596
rect 31276 43540 31332 43550
rect 31276 43446 31332 43484
rect 30716 41858 30772 41870
rect 30716 41806 30718 41858
rect 30770 41806 30772 41858
rect 30716 40964 30772 41806
rect 31164 41860 31220 41870
rect 31164 41766 31220 41804
rect 30716 40180 30772 40908
rect 31724 40292 31780 45052
rect 32284 44996 32340 49200
rect 33180 46116 33236 46126
rect 33180 46022 33236 46060
rect 33628 46116 33684 49200
rect 33628 46050 33684 46060
rect 32284 44930 32340 44940
rect 33068 45892 33124 45902
rect 32732 44210 32788 44222
rect 32732 44158 32734 44210
rect 32786 44158 32788 44210
rect 31724 40226 31780 40236
rect 32508 41860 32564 41870
rect 32508 40290 32564 41804
rect 32732 41412 32788 44158
rect 33068 44210 33124 45836
rect 34972 45332 35028 49200
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35980 45892 36036 45902
rect 35980 45798 36036 45836
rect 34972 45266 35028 45276
rect 34412 45108 34468 45118
rect 33292 44996 33348 45006
rect 33292 44902 33348 44940
rect 33068 44158 33070 44210
rect 33122 44158 33124 44210
rect 33068 44146 33124 44158
rect 33404 44212 33460 44222
rect 33404 44118 33460 44156
rect 33740 44212 33796 44222
rect 33740 44118 33796 44156
rect 34076 44210 34132 44222
rect 34076 44158 34078 44210
rect 34130 44158 34132 44210
rect 33404 43764 33460 43774
rect 33404 43650 33460 43708
rect 33404 43598 33406 43650
rect 33458 43598 33460 43650
rect 33404 43586 33460 43598
rect 33180 43540 33236 43550
rect 33180 43446 33236 43484
rect 32732 41346 32788 41356
rect 32508 40238 32510 40290
rect 32562 40238 32564 40290
rect 30716 40114 30772 40124
rect 31500 40180 31556 40190
rect 30828 39956 30884 39966
rect 30828 39060 30884 39900
rect 30828 38948 30884 39004
rect 30940 38948 30996 38958
rect 30828 38946 30996 38948
rect 30828 38894 30942 38946
rect 30994 38894 30996 38946
rect 30828 38892 30996 38894
rect 30716 38724 30772 38762
rect 30716 38658 30772 38668
rect 30828 35364 30884 38892
rect 30940 38882 30996 38892
rect 31500 38948 31556 40124
rect 32284 39844 32340 39854
rect 32284 39732 32340 39788
rect 32284 39730 32452 39732
rect 32284 39678 32286 39730
rect 32338 39678 32452 39730
rect 32284 39676 32452 39678
rect 32284 39666 32340 39676
rect 32060 38948 32116 38958
rect 31500 38946 32116 38948
rect 31500 38894 31502 38946
rect 31554 38894 32062 38946
rect 32114 38894 32116 38946
rect 31500 38892 32116 38894
rect 31500 38882 31556 38892
rect 32060 38882 32116 38892
rect 32396 38668 32452 39676
rect 32508 39620 32564 40238
rect 32732 39620 32788 39630
rect 32508 39564 32732 39620
rect 32508 39060 32564 39070
rect 32508 38966 32564 39004
rect 32396 38612 32564 38668
rect 32508 37492 32564 38612
rect 32508 37398 32564 37436
rect 32620 36596 32676 39564
rect 32732 39526 32788 39564
rect 33404 39506 33460 39518
rect 33404 39454 33406 39506
rect 33458 39454 33460 39506
rect 33404 39172 33460 39454
rect 33404 39106 33460 39116
rect 33964 39060 34020 39070
rect 34076 39060 34132 44158
rect 34412 44210 34468 45052
rect 35196 45108 35252 45118
rect 35196 45014 35252 45052
rect 35980 45106 36036 45118
rect 35980 45054 35982 45106
rect 36034 45054 36036 45106
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35420 44324 35476 44334
rect 35644 44324 35700 44334
rect 35420 44322 35588 44324
rect 35420 44270 35422 44322
rect 35474 44270 35588 44322
rect 35420 44268 35588 44270
rect 35420 44258 35476 44268
rect 34412 44158 34414 44210
rect 34466 44158 34468 44210
rect 34412 44146 34468 44158
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35532 41524 35588 44268
rect 35644 44210 35700 44268
rect 35644 44158 35646 44210
rect 35698 44158 35700 44210
rect 35644 44146 35700 44158
rect 35980 43764 36036 45054
rect 36316 44548 36372 49200
rect 36988 46116 37044 46126
rect 36988 46022 37044 46060
rect 37660 46116 37716 49200
rect 37660 46050 37716 46060
rect 36988 45332 37044 45342
rect 36988 45238 37044 45276
rect 36316 44482 36372 44492
rect 37996 44548 38052 44558
rect 37996 44454 38052 44492
rect 39004 44548 39060 49200
rect 39788 45890 39844 45902
rect 39788 45838 39790 45890
rect 39842 45838 39844 45890
rect 39788 45556 39844 45838
rect 39788 45490 39844 45500
rect 40348 45332 40404 49200
rect 40796 46116 40852 46126
rect 40796 46022 40852 46060
rect 41692 46116 41748 49200
rect 41692 46050 41748 46060
rect 40348 45266 40404 45276
rect 41916 45332 41972 45342
rect 41916 45238 41972 45276
rect 43036 45332 43092 49200
rect 43036 45266 43092 45276
rect 43932 45890 43988 45902
rect 43932 45838 43934 45890
rect 43986 45838 43988 45890
rect 41020 45106 41076 45118
rect 43820 45108 43876 45118
rect 41020 45054 41022 45106
rect 41074 45054 41076 45106
rect 39004 44482 39060 44492
rect 40908 44548 40964 44558
rect 40908 44454 40964 44492
rect 36988 44324 37044 44334
rect 36988 44230 37044 44268
rect 39900 44322 39956 44334
rect 39900 44270 39902 44322
rect 39954 44270 39956 44322
rect 39900 44212 39956 44270
rect 39900 44146 39956 44156
rect 35980 43698 36036 43708
rect 37324 43540 37380 43550
rect 35532 41468 35812 41524
rect 33964 39058 34132 39060
rect 33964 39006 33966 39058
rect 34018 39006 34132 39058
rect 33964 39004 34132 39006
rect 34188 40292 34244 40302
rect 33964 38994 34020 39004
rect 33292 38724 33348 38762
rect 33292 38612 33460 38668
rect 33180 37492 33236 37502
rect 33236 37436 33348 37492
rect 33180 37426 33236 37436
rect 33292 37378 33348 37436
rect 33292 37326 33294 37378
rect 33346 37326 33348 37378
rect 33292 37314 33348 37326
rect 32620 36594 33124 36596
rect 32620 36542 32622 36594
rect 32674 36542 33124 36594
rect 32620 36540 33124 36542
rect 32620 36530 32676 36540
rect 32172 36260 32228 36270
rect 32172 35810 32228 36204
rect 32172 35758 32174 35810
rect 32226 35758 32228 35810
rect 32172 35746 32228 35758
rect 32396 35810 32452 35822
rect 32396 35758 32398 35810
rect 32450 35758 32452 35810
rect 31836 35588 31892 35598
rect 32396 35588 32452 35758
rect 31836 35586 32452 35588
rect 31836 35534 31838 35586
rect 31890 35534 32452 35586
rect 31836 35532 32452 35534
rect 32508 35588 32564 35598
rect 31836 35522 31892 35532
rect 30604 35086 30606 35138
rect 30658 35086 30660 35138
rect 30604 35074 30660 35086
rect 30716 35308 30884 35364
rect 30268 35028 30324 35066
rect 30268 34962 30324 34972
rect 29820 33346 30212 33348
rect 29820 33294 30158 33346
rect 30210 33294 30212 33346
rect 29820 33292 30212 33294
rect 29708 33236 29764 33246
rect 29708 33142 29764 33180
rect 29708 32450 29764 32462
rect 29708 32398 29710 32450
rect 29762 32398 29764 32450
rect 29708 32116 29764 32398
rect 29820 32338 29876 33292
rect 30156 33282 30212 33292
rect 30268 34804 30324 34814
rect 29820 32286 29822 32338
rect 29874 32286 29876 32338
rect 29820 32274 29876 32286
rect 29708 32050 29764 32060
rect 30156 30210 30212 30222
rect 30156 30158 30158 30210
rect 30210 30158 30212 30210
rect 29708 28644 29764 28654
rect 29708 28530 29764 28588
rect 29708 28478 29710 28530
rect 29762 28478 29764 28530
rect 29708 28466 29764 28478
rect 29932 27748 29988 27758
rect 29932 27654 29988 27692
rect 30156 27524 30212 30158
rect 30268 27860 30324 34748
rect 30380 34130 30436 34142
rect 30380 34078 30382 34130
rect 30434 34078 30436 34130
rect 30380 33908 30436 34078
rect 30604 33908 30660 33918
rect 30380 33906 30660 33908
rect 30380 33854 30606 33906
rect 30658 33854 30660 33906
rect 30380 33852 30660 33854
rect 30604 33842 30660 33852
rect 30380 33236 30436 33246
rect 30380 33142 30436 33180
rect 30716 31556 30772 35308
rect 30828 35140 30884 35150
rect 30828 31892 30884 35084
rect 30940 34018 30996 34030
rect 30940 33966 30942 34018
rect 30994 33966 30996 34018
rect 30940 33906 30996 33966
rect 30940 33854 30942 33906
rect 30994 33854 30996 33906
rect 30940 32004 30996 33854
rect 30940 31948 31332 32004
rect 30828 31890 31220 31892
rect 30828 31838 30830 31890
rect 30882 31838 31220 31890
rect 30828 31836 31220 31838
rect 30828 31826 30884 31836
rect 31164 31778 31220 31836
rect 31164 31726 31166 31778
rect 31218 31726 31220 31778
rect 31164 31714 31220 31726
rect 30716 31500 30884 31556
rect 30380 31108 30436 31118
rect 30380 30212 30436 31052
rect 30380 30210 30548 30212
rect 30380 30158 30382 30210
rect 30434 30158 30548 30210
rect 30380 30156 30548 30158
rect 30380 30146 30436 30156
rect 30492 29314 30548 30156
rect 30716 30100 30772 30110
rect 30716 30006 30772 30044
rect 30492 29262 30494 29314
rect 30546 29262 30548 29314
rect 30492 29250 30548 29262
rect 30268 27794 30324 27804
rect 30156 26908 30212 27468
rect 30828 26908 30884 31500
rect 31164 30212 31220 30222
rect 31276 30212 31332 31948
rect 30940 30156 31164 30212
rect 31220 30156 31332 30212
rect 31836 30324 31892 30334
rect 31836 30210 31892 30268
rect 31836 30158 31838 30210
rect 31890 30158 31892 30210
rect 30940 29652 30996 30156
rect 31164 30118 31220 30156
rect 31836 30146 31892 30158
rect 30940 29558 30996 29596
rect 31276 29540 31332 29550
rect 31276 28084 31332 29484
rect 31948 28420 32004 35532
rect 32508 35494 32564 35532
rect 32732 35028 32788 36540
rect 33068 35698 33124 36540
rect 33068 35646 33070 35698
rect 33122 35646 33124 35698
rect 33068 35634 33124 35646
rect 32732 34934 32788 34972
rect 33404 32788 33460 38612
rect 34188 37492 34244 40236
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34972 39844 35028 39854
rect 34524 38948 34580 38958
rect 34300 38724 34356 38762
rect 34524 38668 34580 38892
rect 34972 38946 35028 39788
rect 35532 39844 35588 39854
rect 35532 39730 35588 39788
rect 35532 39678 35534 39730
rect 35586 39678 35588 39730
rect 35532 39060 35588 39678
rect 35644 39060 35700 39070
rect 35532 39058 35700 39060
rect 35532 39006 35646 39058
rect 35698 39006 35700 39058
rect 35532 39004 35700 39006
rect 35644 38994 35700 39004
rect 34972 38894 34974 38946
rect 35026 38894 35028 38946
rect 34972 38882 35028 38894
rect 34300 38658 34356 38668
rect 34412 38612 34580 38668
rect 34300 37492 34356 37502
rect 34188 37490 34356 37492
rect 34188 37438 34302 37490
rect 34354 37438 34356 37490
rect 34188 37436 34356 37438
rect 34300 37426 34356 37436
rect 33740 37380 33796 37390
rect 33740 37044 33796 37324
rect 33964 37156 34020 37166
rect 33964 37062 34020 37100
rect 33740 34580 33796 36988
rect 33852 35588 33908 35598
rect 33852 35494 33908 35532
rect 33740 34524 33908 34580
rect 32284 32732 33460 32788
rect 33516 34020 33572 34030
rect 31948 28354 32004 28364
rect 32172 28532 32228 28542
rect 31276 28082 31556 28084
rect 31276 28030 31278 28082
rect 31330 28030 31556 28082
rect 31276 28028 31556 28030
rect 31276 28018 31332 28028
rect 31500 27970 31556 28028
rect 31500 27918 31502 27970
rect 31554 27918 31556 27970
rect 31500 27906 31556 27918
rect 31612 27972 31668 27982
rect 31836 27972 31892 27982
rect 32172 27972 32228 28476
rect 31612 27970 31780 27972
rect 31612 27918 31614 27970
rect 31666 27918 31780 27970
rect 31612 27916 31780 27918
rect 31612 27906 31668 27916
rect 31724 27412 31780 27916
rect 31836 27970 32228 27972
rect 31836 27918 31838 27970
rect 31890 27918 32174 27970
rect 32226 27918 32228 27970
rect 31836 27916 32228 27918
rect 31836 27906 31892 27916
rect 32172 27906 32228 27916
rect 31612 27356 31780 27412
rect 31836 27748 31892 27758
rect 30156 26852 30436 26908
rect 30828 26852 30996 26908
rect 29708 24610 29764 24622
rect 29708 24558 29710 24610
rect 29762 24558 29764 24610
rect 29708 24052 29764 24558
rect 29820 24052 29876 24062
rect 29708 24050 29876 24052
rect 29708 23998 29822 24050
rect 29874 23998 29876 24050
rect 29708 23996 29876 23998
rect 29820 23986 29876 23996
rect 29596 23886 29598 23938
rect 29650 23886 29652 23938
rect 29596 23828 29652 23886
rect 30380 23940 30436 26852
rect 30492 24724 30548 24734
rect 30492 24630 30548 24668
rect 30828 24052 30884 24062
rect 30492 23940 30548 23950
rect 30716 23940 30772 23950
rect 30380 23938 30548 23940
rect 30380 23886 30494 23938
rect 30546 23886 30548 23938
rect 30380 23884 30548 23886
rect 30492 23874 30548 23884
rect 30604 23938 30772 23940
rect 30604 23886 30718 23938
rect 30770 23886 30772 23938
rect 30604 23884 30772 23886
rect 29596 23762 29652 23772
rect 29932 23828 29988 23838
rect 30268 23828 30324 23838
rect 29932 23826 30324 23828
rect 29932 23774 29934 23826
rect 29986 23774 30270 23826
rect 30322 23774 30324 23826
rect 29932 23772 30324 23774
rect 29932 23548 29988 23772
rect 30268 23762 30324 23772
rect 29820 23492 29988 23548
rect 28812 22978 28868 22988
rect 29708 23044 29764 23054
rect 29708 22950 29764 22988
rect 29596 22370 29652 22382
rect 29596 22318 29598 22370
rect 29650 22318 29652 22370
rect 29596 22148 29652 22318
rect 29820 22148 29876 23492
rect 30268 23266 30324 23278
rect 30268 23214 30270 23266
rect 30322 23214 30324 23266
rect 30268 23044 30324 23214
rect 30268 22978 30324 22988
rect 30380 23044 30436 23054
rect 30604 23044 30660 23884
rect 30716 23874 30772 23884
rect 30828 23938 30884 23996
rect 30828 23886 30830 23938
rect 30882 23886 30884 23938
rect 30828 23874 30884 23886
rect 30940 23380 30996 26852
rect 31612 26292 31668 27356
rect 31836 26908 31892 27692
rect 31948 27188 32004 27198
rect 31948 27094 32004 27132
rect 31612 26226 31668 26236
rect 31724 26852 31892 26908
rect 31612 25396 31668 25406
rect 31164 25394 31668 25396
rect 31164 25342 31614 25394
rect 31666 25342 31668 25394
rect 31164 25340 31668 25342
rect 31052 24724 31108 24734
rect 31052 24630 31108 24668
rect 31052 23716 31108 23726
rect 31164 23716 31220 25340
rect 31612 25330 31668 25340
rect 31500 23940 31556 23950
rect 31500 23846 31556 23884
rect 31052 23714 31220 23716
rect 31052 23662 31054 23714
rect 31106 23662 31220 23714
rect 31052 23660 31220 23662
rect 31052 23650 31108 23660
rect 30380 23042 30660 23044
rect 30380 22990 30382 23042
rect 30434 22990 30660 23042
rect 30380 22988 30660 22990
rect 30716 23324 30996 23380
rect 30380 22978 30436 22988
rect 29596 22082 29652 22092
rect 29708 22146 29876 22148
rect 29708 22094 29822 22146
rect 29874 22094 29876 22146
rect 29708 22092 29876 22094
rect 29372 20804 29428 20814
rect 29372 20710 29428 20748
rect 29708 20634 29764 22092
rect 29820 22082 29876 22092
rect 30044 22930 30100 22942
rect 30044 22878 30046 22930
rect 30098 22878 30100 22930
rect 30044 22148 30100 22878
rect 30044 22082 30100 22092
rect 30044 21924 30100 21934
rect 29932 20804 29988 20814
rect 29932 20710 29988 20748
rect 29596 20580 29652 20590
rect 28588 20578 29652 20580
rect 28588 20526 28590 20578
rect 28642 20526 29598 20578
rect 29650 20526 29652 20578
rect 28588 20524 29652 20526
rect 28588 18228 28644 20524
rect 29596 20514 29652 20524
rect 29708 20582 29710 20634
rect 29762 20582 29764 20634
rect 29708 19236 29764 20582
rect 29708 19170 29764 19180
rect 29260 19010 29316 19022
rect 29260 18958 29262 19010
rect 29314 18958 29316 19010
rect 29260 18900 29316 18958
rect 28700 18844 29652 18900
rect 28700 18450 28756 18844
rect 29372 18562 29428 18574
rect 29372 18510 29374 18562
rect 29426 18510 29428 18562
rect 28700 18398 28702 18450
rect 28754 18398 28756 18450
rect 28700 18386 28756 18398
rect 29036 18450 29092 18462
rect 29036 18398 29038 18450
rect 29090 18398 29092 18450
rect 28588 18172 28756 18228
rect 28588 17444 28644 17454
rect 28588 17350 28644 17388
rect 28588 15316 28644 15326
rect 28588 15222 28644 15260
rect 28364 15092 28532 15148
rect 28364 14644 28420 15092
rect 28028 14478 28030 14530
rect 28082 14478 28084 14530
rect 28028 14466 28084 14478
rect 28140 14588 28420 14644
rect 27916 14252 28084 14308
rect 27916 13972 27972 13982
rect 27804 13970 27972 13972
rect 27804 13918 27918 13970
rect 27970 13918 27972 13970
rect 27804 13916 27972 13918
rect 27916 13860 27972 13916
rect 27916 13794 27972 13804
rect 28028 13858 28084 14252
rect 28028 13806 28030 13858
rect 28082 13806 28084 13858
rect 28028 13794 28084 13806
rect 27692 13748 27748 13758
rect 27580 13746 27748 13748
rect 27580 13694 27694 13746
rect 27746 13694 27748 13746
rect 27580 13692 27748 13694
rect 27468 12738 27524 12750
rect 27468 12686 27470 12738
rect 27522 12686 27524 12738
rect 27468 12290 27524 12686
rect 27468 12238 27470 12290
rect 27522 12238 27524 12290
rect 27468 12226 27524 12238
rect 27580 12180 27636 13692
rect 27692 13682 27748 13692
rect 27804 13412 27860 13422
rect 27804 12962 27860 13356
rect 28140 12964 28196 14588
rect 27804 12910 27806 12962
rect 27858 12910 27860 12962
rect 27804 12898 27860 12910
rect 27916 12908 28196 12964
rect 28364 14418 28420 14430
rect 28364 14366 28366 14418
rect 28418 14366 28420 14418
rect 27692 12852 27748 12862
rect 27692 12740 27748 12796
rect 27916 12740 27972 12908
rect 27692 12738 27972 12740
rect 27692 12686 27694 12738
rect 27746 12686 27972 12738
rect 27692 12684 27972 12686
rect 27692 12674 27748 12684
rect 27692 12404 27748 12414
rect 27692 12402 28196 12404
rect 27692 12350 27694 12402
rect 27746 12350 28196 12402
rect 27692 12348 28196 12350
rect 27692 12338 27748 12348
rect 27692 12180 27748 12190
rect 27580 12178 27748 12180
rect 27580 12126 27694 12178
rect 27746 12126 27748 12178
rect 27580 12124 27748 12126
rect 27356 12114 27412 12124
rect 27692 12114 27748 12124
rect 27916 12180 27972 12190
rect 27916 12086 27972 12124
rect 28140 11954 28196 12348
rect 28140 11902 28142 11954
rect 28194 11902 28196 11954
rect 28140 11890 28196 11902
rect 27244 10770 27300 10780
rect 26908 9986 26964 9996
rect 26684 8930 26740 8942
rect 26684 8878 26686 8930
rect 26738 8878 26740 8930
rect 26684 8428 26740 8878
rect 27132 8932 27188 8942
rect 27132 8838 27188 8876
rect 28364 8428 28420 14366
rect 28588 14308 28644 14318
rect 28476 13860 28532 13870
rect 28476 13766 28532 13804
rect 28588 13076 28644 14252
rect 28588 12982 28644 13020
rect 28588 12180 28644 12190
rect 28588 12086 28644 12124
rect 28476 11954 28532 11966
rect 28476 11902 28478 11954
rect 28530 11902 28532 11954
rect 28476 10722 28532 11902
rect 28476 10670 28478 10722
rect 28530 10670 28532 10722
rect 28476 10658 28532 10670
rect 26684 8372 27188 8428
rect 26348 8166 26404 8204
rect 27132 4338 27188 8372
rect 28252 8372 28420 8428
rect 28252 6020 28308 8372
rect 28700 6692 28756 18172
rect 29036 18116 29092 18398
rect 29036 18050 29092 18060
rect 29372 17556 29428 18510
rect 29372 17490 29428 17500
rect 29484 17666 29540 17678
rect 29484 17614 29486 17666
rect 29538 17614 29540 17666
rect 29148 17108 29204 17118
rect 29484 17108 29540 17614
rect 29204 17052 29540 17108
rect 29148 17014 29204 17052
rect 29596 16212 29652 18844
rect 30044 18452 30100 21868
rect 30716 21028 30772 23324
rect 30492 20972 30772 21028
rect 30828 23156 30884 23166
rect 30156 20692 30212 20702
rect 30156 20598 30212 20636
rect 30380 20690 30436 20702
rect 30380 20638 30382 20690
rect 30434 20638 30436 20690
rect 30380 20244 30436 20638
rect 30492 20468 30548 20972
rect 30828 20916 30884 23100
rect 31724 21812 31780 26852
rect 31724 21746 31780 21756
rect 32060 21588 32116 21598
rect 30940 20916 30996 20926
rect 30828 20914 30996 20916
rect 30828 20862 30942 20914
rect 30994 20862 30996 20914
rect 30828 20860 30996 20862
rect 30940 20850 30996 20860
rect 30604 20692 30660 20702
rect 30604 20690 30884 20692
rect 30604 20638 30606 20690
rect 30658 20638 30884 20690
rect 30604 20636 30884 20638
rect 30604 20626 30660 20636
rect 30492 20412 30660 20468
rect 30492 20244 30548 20254
rect 30380 20242 30548 20244
rect 30380 20190 30494 20242
rect 30546 20190 30548 20242
rect 30380 20188 30548 20190
rect 30492 20178 30548 20188
rect 30268 20132 30324 20142
rect 30268 19906 30324 20076
rect 30268 19854 30270 19906
rect 30322 19854 30324 19906
rect 30268 19796 30324 19854
rect 30268 19730 30324 19740
rect 30604 19460 30660 20412
rect 30828 20244 30884 20636
rect 30828 20178 30884 20188
rect 31836 20244 31892 20254
rect 30716 20132 30772 20142
rect 30716 20038 30772 20076
rect 31836 20130 31892 20188
rect 31836 20078 31838 20130
rect 31890 20078 31892 20130
rect 30492 19404 30660 19460
rect 30828 20018 30884 20030
rect 30828 19966 30830 20018
rect 30882 19966 30884 20018
rect 30828 19796 30884 19966
rect 30492 19012 30548 19404
rect 30604 19236 30660 19246
rect 30604 19142 30660 19180
rect 30716 19012 30772 19022
rect 30492 18956 30660 19012
rect 30492 18452 30548 18462
rect 29932 18396 30492 18452
rect 29820 18338 29876 18350
rect 29820 18286 29822 18338
rect 29874 18286 29876 18338
rect 29820 18116 29876 18286
rect 29820 18050 29876 18060
rect 29932 17666 29988 18396
rect 30492 18358 30548 18396
rect 29932 17614 29934 17666
rect 29986 17614 29988 17666
rect 29932 17602 29988 17614
rect 30156 17890 30212 17902
rect 30156 17838 30158 17890
rect 30210 17838 30212 17890
rect 30156 16324 30212 17838
rect 30604 17780 30660 18956
rect 30716 18918 30772 18956
rect 30492 17724 30660 17780
rect 30380 17556 30436 17566
rect 30380 17106 30436 17500
rect 30492 17220 30548 17724
rect 30604 17554 30660 17566
rect 30604 17502 30606 17554
rect 30658 17502 30660 17554
rect 30604 17444 30660 17502
rect 30716 17556 30772 17566
rect 30716 17462 30772 17500
rect 30604 17378 30660 17388
rect 30492 17164 30660 17220
rect 30380 17054 30382 17106
rect 30434 17054 30436 17106
rect 30380 17042 30436 17054
rect 30156 16258 30212 16268
rect 29596 16146 29652 16156
rect 29932 15764 29988 15774
rect 29932 15540 29988 15708
rect 30268 15540 30324 15550
rect 29932 15538 30268 15540
rect 29932 15486 29934 15538
rect 29986 15486 30268 15538
rect 29932 15484 30268 15486
rect 29932 15474 29988 15484
rect 30268 15446 30324 15484
rect 30156 15314 30212 15326
rect 30156 15262 30158 15314
rect 30210 15262 30212 15314
rect 29260 15204 29316 15214
rect 28924 14532 28980 14542
rect 28924 13972 28980 14476
rect 28924 13878 28980 13916
rect 29260 12962 29316 15148
rect 30156 15204 30212 15262
rect 30156 15138 30212 15148
rect 30492 15314 30548 15326
rect 30492 15262 30494 15314
rect 30546 15262 30548 15314
rect 30156 14532 30212 14542
rect 30156 14438 30212 14476
rect 29372 13972 29428 13982
rect 29372 13970 29876 13972
rect 29372 13918 29374 13970
rect 29426 13918 29876 13970
rect 29372 13916 29876 13918
rect 29372 13906 29428 13916
rect 29820 13858 29876 13916
rect 29820 13806 29822 13858
rect 29874 13806 29876 13858
rect 29708 13746 29764 13758
rect 29708 13694 29710 13746
rect 29762 13694 29764 13746
rect 29708 13524 29764 13694
rect 29820 13636 29876 13806
rect 30044 13860 30100 13870
rect 30268 13860 30324 13870
rect 30044 13858 30324 13860
rect 30044 13806 30046 13858
rect 30098 13806 30270 13858
rect 30322 13806 30324 13858
rect 30044 13804 30324 13806
rect 30044 13794 30100 13804
rect 30268 13794 30324 13804
rect 30492 13746 30548 15262
rect 30492 13694 30494 13746
rect 30546 13694 30548 13746
rect 30492 13682 30548 13694
rect 29820 13580 30212 13636
rect 29764 13468 30100 13524
rect 29708 13458 29764 13468
rect 29260 12910 29262 12962
rect 29314 12910 29316 12962
rect 29260 12898 29316 12910
rect 29372 13076 29428 13086
rect 29372 12850 29428 13020
rect 30044 12964 30100 13468
rect 30044 12870 30100 12908
rect 29372 12798 29374 12850
rect 29426 12798 29428 12850
rect 29372 12786 29428 12798
rect 29596 12738 29652 12750
rect 29596 12686 29598 12738
rect 29650 12686 29652 12738
rect 29260 12180 29316 12190
rect 29260 12086 29316 12124
rect 29596 12178 29652 12686
rect 29708 12738 29764 12750
rect 29708 12686 29710 12738
rect 29762 12686 29764 12738
rect 29708 12292 29764 12686
rect 29932 12740 29988 12750
rect 29932 12738 30100 12740
rect 29932 12686 29934 12738
rect 29986 12686 30100 12738
rect 29932 12684 30100 12686
rect 29932 12674 29988 12684
rect 30044 12628 30100 12684
rect 29820 12292 29876 12302
rect 29708 12290 29876 12292
rect 29708 12238 29822 12290
rect 29874 12238 29876 12290
rect 29708 12236 29876 12238
rect 29820 12226 29876 12236
rect 29596 12126 29598 12178
rect 29650 12126 29652 12178
rect 29596 12114 29652 12126
rect 29708 12068 29764 12078
rect 29708 12066 29988 12068
rect 29708 12014 29710 12066
rect 29762 12014 29988 12066
rect 29708 12012 29988 12014
rect 29708 12002 29764 12012
rect 29148 11732 29204 11742
rect 29148 10610 29204 11676
rect 29148 10558 29150 10610
rect 29202 10558 29204 10610
rect 29148 10500 29204 10558
rect 29148 9826 29204 10444
rect 29708 10500 29764 10510
rect 29708 10406 29764 10444
rect 29932 9938 29988 12012
rect 30044 11732 30100 12572
rect 30156 11956 30212 13580
rect 30380 13634 30436 13646
rect 30380 13582 30382 13634
rect 30434 13582 30436 13634
rect 30380 13076 30436 13582
rect 30604 13300 30660 17164
rect 30828 16994 30884 19740
rect 31724 19796 31780 19806
rect 31276 19122 31332 19134
rect 31276 19070 31278 19122
rect 31330 19070 31332 19122
rect 30940 19012 30996 19022
rect 31276 19012 31332 19070
rect 31724 19122 31780 19740
rect 31724 19070 31726 19122
rect 31778 19070 31780 19122
rect 31724 19058 31780 19070
rect 31388 19012 31444 19022
rect 30940 19010 31220 19012
rect 30940 18958 30942 19010
rect 30994 18958 31220 19010
rect 30940 18956 31220 18958
rect 31276 18956 31388 19012
rect 30940 18946 30996 18956
rect 31164 17668 31220 18956
rect 31388 18946 31444 18956
rect 31836 18564 31892 20078
rect 32060 20018 32116 21532
rect 32060 19966 32062 20018
rect 32114 19966 32116 20018
rect 32060 19954 32116 19966
rect 31948 19908 32004 19918
rect 31948 19234 32004 19852
rect 31948 19182 31950 19234
rect 32002 19182 32004 19234
rect 31948 19170 32004 19182
rect 32172 19348 32228 19358
rect 31836 18508 32004 18564
rect 31388 18340 31444 18350
rect 31388 18246 31444 18284
rect 31836 18340 31892 18350
rect 31836 18246 31892 18284
rect 31276 17668 31332 17678
rect 31612 17668 31668 17678
rect 31164 17666 31332 17668
rect 31164 17614 31278 17666
rect 31330 17614 31332 17666
rect 31164 17612 31332 17614
rect 31276 17602 31332 17612
rect 31388 17666 31668 17668
rect 31388 17614 31614 17666
rect 31666 17614 31668 17666
rect 31388 17612 31668 17614
rect 30940 17444 30996 17454
rect 30940 17442 31108 17444
rect 30940 17390 30942 17442
rect 30994 17390 31108 17442
rect 30940 17388 31108 17390
rect 30940 17378 30996 17388
rect 30940 17220 30996 17230
rect 30940 17106 30996 17164
rect 30940 17054 30942 17106
rect 30994 17054 30996 17106
rect 30940 17042 30996 17054
rect 30828 16942 30830 16994
rect 30882 16942 30884 16994
rect 30828 16660 30884 16942
rect 30828 16604 30996 16660
rect 30940 15988 30996 16604
rect 30940 15922 30996 15932
rect 30716 15876 30772 15886
rect 30716 14308 30772 15820
rect 31052 15148 31108 17388
rect 31388 17220 31444 17612
rect 31612 17602 31668 17612
rect 31948 17556 32004 18508
rect 32172 18450 32228 19292
rect 32172 18398 32174 18450
rect 32226 18398 32228 18450
rect 32172 18386 32228 18398
rect 31836 17554 32004 17556
rect 31836 17502 31950 17554
rect 32002 17502 32004 17554
rect 31836 17500 32004 17502
rect 31612 17442 31668 17454
rect 31612 17390 31614 17442
rect 31666 17390 31668 17442
rect 31164 17164 31444 17220
rect 31500 17220 31556 17230
rect 31164 17106 31220 17164
rect 31164 17054 31166 17106
rect 31218 17054 31220 17106
rect 31164 17042 31220 17054
rect 31500 17106 31556 17164
rect 31500 17054 31502 17106
rect 31554 17054 31556 17106
rect 31500 17042 31556 17054
rect 31612 16660 31668 17390
rect 31612 16594 31668 16604
rect 31724 16996 31780 17006
rect 31164 16100 31220 16110
rect 31164 15876 31220 16044
rect 31500 16100 31556 16110
rect 31388 15988 31444 15998
rect 31388 15894 31444 15932
rect 31500 15986 31556 16044
rect 31724 16098 31780 16940
rect 31724 16046 31726 16098
rect 31778 16046 31780 16098
rect 31724 16034 31780 16046
rect 31500 15934 31502 15986
rect 31554 15934 31556 15986
rect 31500 15922 31556 15934
rect 31836 15876 31892 17500
rect 31948 17490 32004 17500
rect 32060 16212 32116 16222
rect 32060 16098 32116 16156
rect 32060 16046 32062 16098
rect 32114 16046 32116 16098
rect 32060 16034 32116 16046
rect 31164 15782 31220 15820
rect 31612 15820 31892 15876
rect 31052 15092 31444 15148
rect 30716 14242 30772 14252
rect 30828 13860 30884 13870
rect 30828 13766 30884 13804
rect 31052 13748 31108 13758
rect 30604 13234 30660 13244
rect 30940 13746 31108 13748
rect 30940 13694 31054 13746
rect 31106 13694 31108 13746
rect 30940 13692 31108 13694
rect 30380 13020 30660 13076
rect 30268 12964 30324 12974
rect 30268 12852 30324 12908
rect 30380 12852 30436 12862
rect 30268 12850 30436 12852
rect 30268 12798 30382 12850
rect 30434 12798 30436 12850
rect 30268 12796 30436 12798
rect 30380 12786 30436 12796
rect 30492 12740 30548 12750
rect 30492 12646 30548 12684
rect 30380 12180 30436 12190
rect 30380 12086 30436 12124
rect 30156 11890 30212 11900
rect 30044 11676 30324 11732
rect 29932 9886 29934 9938
rect 29986 9886 29988 9938
rect 29932 9874 29988 9886
rect 29148 9774 29150 9826
rect 29202 9774 29204 9826
rect 29148 9762 29204 9774
rect 30268 9604 30324 11676
rect 30604 11508 30660 13020
rect 30716 12964 30772 12974
rect 30940 12964 30996 13692
rect 31052 13682 31108 13692
rect 31388 13746 31444 15092
rect 31388 13694 31390 13746
rect 31442 13694 31444 13746
rect 31388 13682 31444 13694
rect 31612 13860 31668 15820
rect 31724 15540 31780 15550
rect 31948 15540 32004 15550
rect 31780 15538 32004 15540
rect 31780 15486 31950 15538
rect 32002 15486 32004 15538
rect 31780 15484 32004 15486
rect 31724 15446 31780 15484
rect 31948 15474 32004 15484
rect 31612 13746 31668 13804
rect 31612 13694 31614 13746
rect 31666 13694 31668 13746
rect 31612 13682 31668 13694
rect 32060 14418 32116 14430
rect 32060 14366 32062 14418
rect 32114 14366 32116 14418
rect 31276 13634 31332 13646
rect 31276 13582 31278 13634
rect 31330 13582 31332 13634
rect 30716 12962 30996 12964
rect 30716 12910 30718 12962
rect 30770 12910 30996 12962
rect 30716 12908 30996 12910
rect 31052 13300 31108 13310
rect 30716 12898 30772 12908
rect 31052 12738 31108 13244
rect 31276 13076 31332 13582
rect 31276 13010 31332 13020
rect 31388 13524 31444 13534
rect 31052 12686 31054 12738
rect 31106 12686 31108 12738
rect 31052 12628 31108 12686
rect 31052 12562 31108 12572
rect 30604 11442 30660 11452
rect 30940 11732 30996 11742
rect 30940 11394 30996 11676
rect 30940 11342 30942 11394
rect 30994 11342 30996 11394
rect 30940 11330 30996 11342
rect 30268 9538 30324 9548
rect 31388 8428 31444 13468
rect 32060 12962 32116 14366
rect 32060 12910 32062 12962
rect 32114 12910 32116 12962
rect 31500 12740 31556 12750
rect 31500 12646 31556 12684
rect 31612 12068 31668 12078
rect 31612 12066 31892 12068
rect 31612 12014 31614 12066
rect 31666 12014 31892 12066
rect 31612 12012 31892 12014
rect 31612 12002 31668 12012
rect 31836 11844 31892 12012
rect 31948 11844 32004 11854
rect 32060 11844 32116 12910
rect 31836 11788 31948 11844
rect 32004 11788 32116 11844
rect 31948 11750 32004 11788
rect 31612 11508 31668 11518
rect 31668 11452 31780 11508
rect 31612 11442 31668 11452
rect 31724 11394 31780 11452
rect 31724 11342 31726 11394
rect 31778 11342 31780 11394
rect 31724 11330 31780 11342
rect 32172 9604 32228 9614
rect 32172 9510 32228 9548
rect 32284 9156 32340 32732
rect 33516 32228 33572 33964
rect 33516 32172 33796 32228
rect 33628 32004 33684 32014
rect 33516 31948 33628 32004
rect 32732 31220 32788 31230
rect 32396 28420 32452 28430
rect 32396 28082 32452 28364
rect 32396 28030 32398 28082
rect 32450 28030 32452 28082
rect 32396 27188 32452 28030
rect 32508 27748 32564 27758
rect 32508 27654 32564 27692
rect 32396 27122 32452 27132
rect 32732 25732 32788 31164
rect 33068 30212 33124 30222
rect 33068 27858 33124 30156
rect 33516 29650 33572 31948
rect 33628 31938 33684 31948
rect 33516 29598 33518 29650
rect 33570 29598 33572 29650
rect 33516 29586 33572 29598
rect 33628 31668 33684 31678
rect 33180 29426 33236 29438
rect 33180 29374 33182 29426
rect 33234 29374 33236 29426
rect 33180 29204 33236 29374
rect 33180 29138 33236 29148
rect 33628 28084 33684 31612
rect 33740 31220 33796 32172
rect 33852 32116 33908 34524
rect 34188 33570 34244 33582
rect 34188 33518 34190 33570
rect 34242 33518 34244 33570
rect 34076 33236 34132 33246
rect 33852 32050 33908 32060
rect 33964 33180 34076 33236
rect 33740 31126 33796 31164
rect 33852 31780 33908 31790
rect 33852 31108 33908 31724
rect 33852 30324 33908 31052
rect 33964 30772 34020 33180
rect 34076 33170 34132 33180
rect 34188 31668 34244 33518
rect 34412 32788 34468 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34860 37380 34916 37390
rect 34860 37286 34916 37324
rect 35420 37156 35476 37166
rect 35420 37062 35476 37100
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34748 36260 34804 36270
rect 34524 35140 34580 35150
rect 34524 33570 34580 35084
rect 34748 35138 34804 36204
rect 34748 35086 34750 35138
rect 34802 35086 34804 35138
rect 34748 35074 34804 35086
rect 35084 35588 35140 35598
rect 35084 34914 35140 35532
rect 35532 35476 35588 35486
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 34862 35086 34914
rect 35138 34862 35140 34914
rect 35084 34850 35140 34862
rect 34860 34692 34916 34702
rect 34524 33518 34526 33570
rect 34578 33518 34580 33570
rect 34524 33458 34580 33518
rect 34524 33406 34526 33458
rect 34578 33406 34580 33458
rect 34524 33012 34580 33406
rect 34524 32946 34580 32956
rect 34636 34690 34916 34692
rect 34636 34638 34862 34690
rect 34914 34638 34916 34690
rect 34636 34636 34916 34638
rect 34412 32722 34468 32732
rect 34524 32676 34580 32686
rect 34412 32452 34468 32462
rect 34524 32452 34580 32620
rect 34412 32450 34580 32452
rect 34412 32398 34414 32450
rect 34466 32398 34580 32450
rect 34412 32396 34580 32398
rect 34412 32386 34468 32396
rect 34188 31602 34244 31612
rect 34412 31666 34468 31678
rect 34412 31614 34414 31666
rect 34466 31614 34468 31666
rect 34076 31556 34132 31566
rect 34076 31106 34132 31500
rect 34188 31220 34244 31230
rect 34188 31126 34244 31164
rect 34076 31054 34078 31106
rect 34130 31054 34132 31106
rect 34076 30996 34132 31054
rect 34076 30930 34132 30940
rect 34188 30772 34244 30782
rect 33964 30770 34244 30772
rect 33964 30718 34190 30770
rect 34242 30718 34244 30770
rect 33964 30716 34244 30718
rect 34188 30706 34244 30716
rect 34188 30548 34244 30558
rect 33964 30324 34020 30334
rect 33852 30322 34020 30324
rect 33852 30270 33966 30322
rect 34018 30270 34020 30322
rect 33852 30268 34020 30270
rect 33964 30258 34020 30268
rect 33628 28018 33684 28028
rect 33068 27806 33070 27858
rect 33122 27806 33124 27858
rect 33068 26908 33124 27806
rect 33852 27748 33908 27758
rect 33852 27654 33908 27692
rect 34188 26908 34244 30492
rect 34412 30322 34468 31614
rect 34412 30270 34414 30322
rect 34466 30270 34468 30322
rect 34412 30212 34468 30270
rect 34412 30146 34468 30156
rect 34524 29988 34580 32396
rect 34412 29932 34580 29988
rect 34412 27972 34468 29932
rect 34636 29540 34692 34636
rect 34860 34626 34916 34636
rect 35532 34354 35588 35420
rect 35532 34302 35534 34354
rect 35586 34302 35588 34354
rect 35532 34290 35588 34302
rect 35196 34132 35252 34142
rect 34972 34130 35252 34132
rect 34972 34078 35198 34130
rect 35250 34078 35252 34130
rect 34972 34076 35252 34078
rect 34972 33570 35028 34076
rect 35196 34066 35252 34076
rect 35532 34130 35588 34142
rect 35532 34078 35534 34130
rect 35586 34078 35588 34130
rect 35532 33908 35588 34078
rect 35532 33842 35588 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34972 33518 34974 33570
rect 35026 33518 35028 33570
rect 34972 33506 35028 33518
rect 35532 33460 35588 33470
rect 35756 33460 35812 41468
rect 35980 39620 36036 39630
rect 35980 39526 36036 39564
rect 36092 38948 36148 38958
rect 36092 38854 36148 38892
rect 36652 38724 36708 38762
rect 36652 38658 36708 38668
rect 35868 37156 35924 37166
rect 35868 35364 35924 37100
rect 36428 35698 36484 35710
rect 36428 35646 36430 35698
rect 36482 35646 36484 35698
rect 35980 35588 36036 35598
rect 35980 35494 36036 35532
rect 35868 35308 36036 35364
rect 35532 33366 35588 33404
rect 35644 33404 35812 33460
rect 35868 34130 35924 34142
rect 35868 34078 35870 34130
rect 35922 34078 35924 34130
rect 35308 33348 35364 33358
rect 35084 33346 35364 33348
rect 35084 33294 35310 33346
rect 35362 33294 35364 33346
rect 35084 33292 35364 33294
rect 34748 33180 34916 33236
rect 34748 32562 34804 33180
rect 34860 33178 34916 33180
rect 34860 33126 34862 33178
rect 34914 33126 34916 33178
rect 34860 33114 34916 33126
rect 34972 33122 35028 33134
rect 34972 33070 34974 33122
rect 35026 33070 35028 33122
rect 34860 33012 34916 33022
rect 34972 33012 35028 33070
rect 34916 32956 35028 33012
rect 34860 32946 34916 32956
rect 35084 32786 35140 33292
rect 35308 33282 35364 33292
rect 35644 32900 35700 33404
rect 35868 33348 35924 34078
rect 35756 33236 35812 33246
rect 35756 33142 35812 33180
rect 35084 32734 35086 32786
rect 35138 32734 35140 32786
rect 35084 32722 35140 32734
rect 35532 32844 35700 32900
rect 34860 32676 34916 32686
rect 34860 32582 34916 32620
rect 35420 32674 35476 32686
rect 35420 32622 35422 32674
rect 35474 32622 35476 32674
rect 34748 32510 34750 32562
rect 34802 32510 34804 32562
rect 34748 32452 34804 32510
rect 35308 32562 35364 32574
rect 35308 32510 35310 32562
rect 35362 32510 35364 32562
rect 35308 32452 35364 32510
rect 34748 32396 35364 32452
rect 34748 32004 34804 32396
rect 35420 32340 35476 32622
rect 35420 32274 35476 32284
rect 35532 32228 35588 32844
rect 35644 32674 35700 32686
rect 35644 32622 35646 32674
rect 35698 32622 35700 32674
rect 35644 32564 35700 32622
rect 35756 32564 35812 32574
rect 35644 32508 35756 32564
rect 35756 32498 35812 32508
rect 35868 32562 35924 33292
rect 35868 32510 35870 32562
rect 35922 32510 35924 32562
rect 35868 32498 35924 32510
rect 35196 32172 35460 32182
rect 35532 32172 35924 32228
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34748 31938 34804 31948
rect 35868 31218 35924 32172
rect 35868 31166 35870 31218
rect 35922 31166 35924 31218
rect 35868 31154 35924 31166
rect 34860 31108 34916 31118
rect 34860 31014 34916 31052
rect 34748 30994 34804 31006
rect 35980 30996 36036 35308
rect 36092 35028 36148 35038
rect 36428 35028 36484 35646
rect 37212 35586 37268 35598
rect 37212 35534 37214 35586
rect 37266 35534 37268 35586
rect 37212 35476 37268 35534
rect 37212 35410 37268 35420
rect 36148 34972 36484 35028
rect 36092 34934 36148 34972
rect 36876 32788 36932 32798
rect 36092 32562 36148 32574
rect 36092 32510 36094 32562
rect 36146 32510 36148 32562
rect 36092 31220 36148 32510
rect 36428 32564 36484 32574
rect 36428 32470 36484 32508
rect 36316 32452 36372 32462
rect 36316 32358 36372 32396
rect 36876 32450 36932 32732
rect 36876 32398 36878 32450
rect 36930 32398 36932 32450
rect 36876 32340 36932 32398
rect 36876 32274 36932 32284
rect 36876 32004 36932 32014
rect 36204 31220 36260 31230
rect 36092 31218 36260 31220
rect 36092 31166 36206 31218
rect 36258 31166 36260 31218
rect 36092 31164 36260 31166
rect 36204 31154 36260 31164
rect 34748 30942 34750 30994
rect 34802 30942 34804 30994
rect 34748 30436 34804 30942
rect 35868 30940 36036 30996
rect 36428 31106 36484 31118
rect 36428 31054 36430 31106
rect 36482 31054 36484 31106
rect 34748 30370 34804 30380
rect 34860 30884 34916 30894
rect 34636 29474 34692 29484
rect 34860 29538 34916 30828
rect 35532 30770 35588 30782
rect 35532 30718 35534 30770
rect 35586 30718 35588 30770
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35532 30324 35588 30718
rect 35532 30258 35588 30268
rect 35308 30098 35364 30110
rect 35532 30100 35588 30110
rect 35308 30046 35310 30098
rect 35362 30046 35364 30098
rect 35084 29988 35140 29998
rect 35308 29988 35364 30046
rect 35084 29986 35364 29988
rect 35084 29934 35086 29986
rect 35138 29934 35364 29986
rect 35084 29932 35364 29934
rect 35420 30098 35588 30100
rect 35420 30046 35534 30098
rect 35586 30046 35588 30098
rect 35420 30044 35588 30046
rect 34860 29486 34862 29538
rect 34914 29486 34916 29538
rect 34860 29474 34916 29486
rect 34972 29538 35028 29550
rect 34972 29486 34974 29538
rect 35026 29486 35028 29538
rect 34412 27906 34468 27916
rect 34524 29314 34580 29326
rect 34524 29262 34526 29314
rect 34578 29262 34580 29314
rect 34524 29204 34580 29262
rect 34972 29204 35028 29486
rect 34524 29148 35028 29204
rect 33068 26852 33572 26908
rect 33180 26178 33236 26190
rect 33180 26126 33182 26178
rect 33234 26126 33236 26178
rect 32508 25676 32788 25732
rect 32844 25844 32900 25854
rect 32396 25620 32452 25630
rect 32396 25506 32452 25564
rect 32396 25454 32398 25506
rect 32450 25454 32452 25506
rect 32396 25442 32452 25454
rect 32508 19124 32564 25676
rect 32844 25618 32900 25788
rect 32844 25566 32846 25618
rect 32898 25566 32900 25618
rect 32844 25554 32900 25566
rect 33180 25282 33236 26126
rect 33180 25230 33182 25282
rect 33234 25230 33236 25282
rect 33180 23044 33236 25230
rect 33292 25620 33348 26852
rect 33516 26786 33572 26796
rect 34076 26852 34244 26908
rect 34524 26908 34580 29148
rect 35084 28980 35140 29932
rect 35420 29764 35476 30044
rect 35532 30034 35588 30044
rect 35756 30100 35812 30110
rect 35756 30006 35812 30044
rect 35196 29708 35476 29764
rect 35196 29650 35252 29708
rect 35196 29598 35198 29650
rect 35250 29598 35252 29650
rect 35196 29586 35252 29598
rect 35420 29540 35476 29550
rect 35476 29484 35588 29540
rect 35420 29474 35476 29484
rect 34972 28924 35140 28980
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34860 28644 34916 28654
rect 34972 28644 35028 28924
rect 34916 28588 35028 28644
rect 35084 28754 35140 28766
rect 35084 28702 35086 28754
rect 35138 28702 35140 28754
rect 34860 28578 34916 28588
rect 34748 28532 34804 28542
rect 34748 28438 34804 28476
rect 34972 28418 35028 28430
rect 34972 28366 34974 28418
rect 35026 28366 35028 28418
rect 34972 27748 35028 28366
rect 34972 27682 35028 27692
rect 35084 27076 35140 28702
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35532 27300 35588 29484
rect 35420 27244 35588 27300
rect 35308 27076 35364 27086
rect 35084 27074 35364 27076
rect 35084 27022 35310 27074
rect 35362 27022 35364 27074
rect 35084 27020 35364 27022
rect 35308 27010 35364 27020
rect 34524 26852 34804 26908
rect 33292 24946 33348 25564
rect 33404 26180 33460 26190
rect 33404 25506 33460 26124
rect 33740 26178 33796 26190
rect 33740 26126 33742 26178
rect 33794 26126 33796 26178
rect 33516 25956 33572 25966
rect 33516 25730 33572 25900
rect 33516 25678 33518 25730
rect 33570 25678 33572 25730
rect 33516 25666 33572 25678
rect 33628 25844 33684 25854
rect 33404 25454 33406 25506
rect 33458 25454 33460 25506
rect 33404 25396 33460 25454
rect 33628 25508 33684 25788
rect 33740 25508 33796 26126
rect 33964 25508 34020 25518
rect 33628 25506 34020 25508
rect 33628 25454 33630 25506
rect 33682 25454 33966 25506
rect 34018 25454 34020 25506
rect 33628 25452 34020 25454
rect 33628 25442 33684 25452
rect 33964 25442 34020 25452
rect 33404 25330 33460 25340
rect 33292 24894 33294 24946
rect 33346 24894 33348 24946
rect 33292 24882 33348 24894
rect 33852 24836 33908 24846
rect 34076 24836 34132 26852
rect 34524 26740 34580 26750
rect 34412 26516 34468 26526
rect 34300 25844 34356 25854
rect 34188 25396 34244 25406
rect 34188 25302 34244 25340
rect 33628 24780 33852 24836
rect 33628 24722 33684 24780
rect 33852 24770 33908 24780
rect 33964 24780 34132 24836
rect 34300 25060 34356 25788
rect 33628 24670 33630 24722
rect 33682 24670 33684 24722
rect 33628 24658 33684 24670
rect 33180 22978 33236 22988
rect 33628 24500 33684 24510
rect 33068 20692 33124 20702
rect 33068 20598 33124 20636
rect 32396 19068 32564 19124
rect 32844 19348 32900 19358
rect 32396 15652 32452 19068
rect 32732 19010 32788 19022
rect 32732 18958 32734 19010
rect 32786 18958 32788 19010
rect 32508 18340 32564 18350
rect 32732 18340 32788 18958
rect 32508 18338 32676 18340
rect 32508 18286 32510 18338
rect 32562 18286 32676 18338
rect 32508 18284 32676 18286
rect 32508 18274 32564 18284
rect 32396 15202 32452 15596
rect 32396 15150 32398 15202
rect 32450 15150 32452 15202
rect 32396 15138 32452 15150
rect 32284 9090 32340 9100
rect 31164 8372 31444 8428
rect 32620 8428 32676 18284
rect 32732 18274 32788 18284
rect 32844 17778 32900 19292
rect 33628 19012 33684 24444
rect 33852 20916 33908 20926
rect 33852 20802 33908 20860
rect 33852 20750 33854 20802
rect 33906 20750 33908 20802
rect 33852 20738 33908 20750
rect 33628 18946 33684 18956
rect 32844 17726 32846 17778
rect 32898 17726 32900 17778
rect 32844 17714 32900 17726
rect 33292 18450 33348 18462
rect 33292 18398 33294 18450
rect 33346 18398 33348 18450
rect 33292 18340 33348 18398
rect 33180 17220 33236 17230
rect 33180 16994 33236 17164
rect 33180 16942 33182 16994
rect 33234 16942 33236 16994
rect 33068 16882 33124 16894
rect 33068 16830 33070 16882
rect 33122 16830 33124 16882
rect 32732 16660 32788 16670
rect 32732 16210 32788 16604
rect 32732 16158 32734 16210
rect 32786 16158 32788 16210
rect 32732 16146 32788 16158
rect 33068 15988 33124 16830
rect 33068 15922 33124 15932
rect 33180 15540 33236 16942
rect 33180 15474 33236 15484
rect 33292 14532 33348 18284
rect 33740 17220 33796 17230
rect 33740 17106 33796 17164
rect 33740 17054 33742 17106
rect 33794 17054 33796 17106
rect 33740 17042 33796 17054
rect 33404 16884 33460 16894
rect 33404 16790 33460 16828
rect 33292 14466 33348 14476
rect 33628 16324 33684 16334
rect 32732 13076 32788 13086
rect 32732 12982 32788 13020
rect 32732 11172 32788 11182
rect 32732 10500 32788 11116
rect 32732 9938 32788 10444
rect 32732 9886 32734 9938
rect 32786 9886 32788 9938
rect 32732 9874 32788 9886
rect 32620 8372 33236 8428
rect 31164 7700 31220 8372
rect 31164 7634 31220 7644
rect 28700 6626 28756 6636
rect 28252 5954 28308 5964
rect 29036 6020 29092 6030
rect 27132 4286 27134 4338
rect 27186 4286 27188 4338
rect 27132 4274 27188 4286
rect 26908 4116 26964 4126
rect 26124 3556 26180 3566
rect 26012 3500 26124 3556
rect 26124 3490 26180 3500
rect 24892 3332 25396 3388
rect 22652 2380 22932 2436
rect 22876 800 22932 2380
rect 24892 800 24948 3332
rect 26908 800 26964 4060
rect 28140 4116 28196 4126
rect 28140 4022 28196 4060
rect 27244 3556 27300 3566
rect 27244 3462 27300 3500
rect 28476 3556 28532 3566
rect 28476 3462 28532 3500
rect 29036 3554 29092 5964
rect 33180 4338 33236 8372
rect 33180 4286 33182 4338
rect 33234 4286 33236 4338
rect 33180 4274 33236 4286
rect 32956 4116 33012 4126
rect 29036 3502 29038 3554
rect 29090 3502 29092 3554
rect 29036 3490 29092 3502
rect 32620 3556 32676 3566
rect 32620 3462 32676 3500
rect 28924 3444 28980 3454
rect 28924 800 28980 3388
rect 30044 3444 30100 3454
rect 30044 3330 30100 3388
rect 30044 3278 30046 3330
rect 30098 3278 30100 3330
rect 30044 3266 30100 3278
rect 30940 3444 30996 3454
rect 30940 800 30996 3388
rect 32956 800 33012 4060
rect 33628 3556 33684 16268
rect 33964 11732 34020 24780
rect 34300 24722 34356 25004
rect 34412 25394 34468 26460
rect 34524 25730 34580 26684
rect 34524 25678 34526 25730
rect 34578 25678 34580 25730
rect 34524 25666 34580 25678
rect 34636 25956 34692 25966
rect 34636 25506 34692 25900
rect 34636 25454 34638 25506
rect 34690 25454 34692 25506
rect 34636 25442 34692 25454
rect 34412 25342 34414 25394
rect 34466 25342 34468 25394
rect 34412 24948 34468 25342
rect 34524 25396 34580 25406
rect 34524 24948 34580 25340
rect 34748 25172 34804 26852
rect 35420 26068 35476 27244
rect 35868 27188 35924 30940
rect 35980 30772 36036 30782
rect 35980 30210 36036 30716
rect 35980 30158 35982 30210
rect 36034 30158 36036 30210
rect 35980 30146 36036 30158
rect 36316 29988 36372 29998
rect 36428 29988 36484 31054
rect 36876 31106 36932 31948
rect 36988 31892 37044 31902
rect 36988 31220 37044 31836
rect 37324 31668 37380 43484
rect 40908 42754 40964 42766
rect 40908 42702 40910 42754
rect 40962 42702 40964 42754
rect 39788 42644 39844 42654
rect 40796 42644 40852 42654
rect 39788 42550 39844 42588
rect 40572 42588 40796 42644
rect 39228 42532 39284 42542
rect 39004 38050 39060 38062
rect 39004 37998 39006 38050
rect 39058 37998 39060 38050
rect 39004 37828 39060 37998
rect 39116 37940 39172 37950
rect 39116 37846 39172 37884
rect 38668 35812 38724 35822
rect 38108 33346 38164 33358
rect 38108 33294 38110 33346
rect 38162 33294 38164 33346
rect 37772 33124 37828 33134
rect 38108 33124 38164 33294
rect 37772 33122 38164 33124
rect 37772 33070 37774 33122
rect 37826 33070 38164 33122
rect 37772 33068 38164 33070
rect 37212 31612 37380 31668
rect 37436 32564 37492 32574
rect 37772 32564 37828 33068
rect 37436 32562 37828 32564
rect 37436 32510 37438 32562
rect 37490 32510 37828 32562
rect 37436 32508 37828 32510
rect 36988 31126 37044 31164
rect 37100 31556 37156 31566
rect 36876 31054 36878 31106
rect 36930 31054 36932 31106
rect 36876 31042 36932 31054
rect 36540 30996 36596 31006
rect 36540 30902 36596 30940
rect 36988 30772 37044 30782
rect 36988 30678 37044 30716
rect 36316 29986 36484 29988
rect 36316 29934 36318 29986
rect 36370 29934 36484 29986
rect 36316 29932 36484 29934
rect 36316 29922 36372 29932
rect 35980 29316 36036 29326
rect 35980 28756 36036 29260
rect 35980 28754 36372 28756
rect 35980 28702 35982 28754
rect 36034 28702 36372 28754
rect 35980 28700 36372 28702
rect 35980 28690 36036 28700
rect 36316 28082 36372 28700
rect 36316 28030 36318 28082
rect 36370 28030 36372 28082
rect 36316 28018 36372 28030
rect 35980 27748 36036 27758
rect 35980 27654 36036 27692
rect 35644 27132 35924 27188
rect 35532 27076 35588 27086
rect 35532 26982 35588 27020
rect 35420 26012 35588 26068
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35084 25620 35140 25630
rect 34972 25508 35028 25518
rect 34860 25396 34916 25406
rect 34860 25302 34916 25340
rect 34748 25116 34916 25172
rect 34636 24948 34692 24958
rect 34524 24946 34692 24948
rect 34524 24894 34638 24946
rect 34690 24894 34692 24946
rect 34524 24892 34692 24894
rect 34412 24882 34468 24892
rect 34636 24882 34692 24892
rect 34748 24836 34804 24846
rect 34748 24724 34804 24780
rect 34300 24670 34302 24722
rect 34354 24670 34356 24722
rect 34300 24658 34356 24670
rect 34524 24668 34804 24724
rect 34860 24834 34916 25116
rect 34972 24946 35028 25452
rect 35084 25506 35140 25564
rect 35084 25454 35086 25506
rect 35138 25454 35140 25506
rect 35084 25442 35140 25454
rect 35308 25508 35364 25518
rect 35532 25508 35588 26012
rect 35308 25506 35588 25508
rect 35308 25454 35310 25506
rect 35362 25454 35588 25506
rect 35308 25452 35588 25454
rect 35308 25442 35364 25452
rect 34972 24894 34974 24946
rect 35026 24894 35028 24946
rect 34972 24882 35028 24894
rect 34860 24782 34862 24834
rect 34914 24782 34916 24834
rect 34076 24612 34132 24622
rect 34076 24518 34132 24556
rect 34412 24276 34468 24286
rect 34076 24164 34132 24174
rect 34076 24050 34132 24108
rect 34076 23998 34078 24050
rect 34130 23998 34132 24050
rect 34076 23986 34132 23998
rect 34412 23548 34468 24220
rect 34300 23492 34468 23548
rect 34188 22148 34244 22158
rect 34188 20802 34244 22092
rect 34188 20750 34190 20802
rect 34242 20750 34244 20802
rect 34188 20738 34244 20750
rect 34300 15148 34356 23492
rect 34412 21812 34468 21822
rect 34412 21718 34468 21756
rect 34524 20804 34580 24668
rect 34860 24612 34916 24782
rect 34860 24546 34916 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21812 35252 21822
rect 35196 21718 35252 21756
rect 34748 21698 34804 21710
rect 34748 21646 34750 21698
rect 34802 21646 34804 21698
rect 34748 21588 34804 21646
rect 34748 21522 34804 21532
rect 35420 21588 35476 21598
rect 35476 21532 35588 21588
rect 35420 21522 35476 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34972 20916 35028 20926
rect 34972 20822 35028 20860
rect 34412 20748 34916 20804
rect 34412 20132 34468 20748
rect 34860 20692 34916 20748
rect 35532 20802 35588 21532
rect 35532 20750 35534 20802
rect 35586 20750 35588 20802
rect 35532 20738 35588 20750
rect 34860 20636 35028 20692
rect 34524 20580 34580 20590
rect 34524 20578 34692 20580
rect 34524 20526 34526 20578
rect 34578 20526 34692 20578
rect 34524 20524 34692 20526
rect 34524 20514 34580 20524
rect 34524 20132 34580 20142
rect 34412 20130 34580 20132
rect 34412 20078 34526 20130
rect 34578 20078 34580 20130
rect 34412 20076 34580 20078
rect 34412 17556 34468 20076
rect 34524 20066 34580 20076
rect 34636 19236 34692 20524
rect 34972 20130 35028 20636
rect 34972 20078 34974 20130
rect 35026 20078 35028 20130
rect 34972 20066 35028 20078
rect 35084 20132 35140 20142
rect 34860 20018 34916 20030
rect 34860 19966 34862 20018
rect 34914 19966 34916 20018
rect 34860 19908 34916 19966
rect 34860 19842 34916 19852
rect 35084 19348 35140 20076
rect 35532 20132 35588 20142
rect 35532 20038 35588 20076
rect 35196 20020 35252 20030
rect 35196 19926 35252 19964
rect 35420 20018 35476 20030
rect 35420 19966 35422 20018
rect 35474 19966 35476 20018
rect 35420 19908 35476 19966
rect 35420 19842 35476 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 19348 35252 19358
rect 35084 19346 35252 19348
rect 35084 19294 35198 19346
rect 35250 19294 35252 19346
rect 35084 19292 35252 19294
rect 35196 19282 35252 19292
rect 34636 19170 34692 19180
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34412 17490 34468 17500
rect 35420 17108 35476 17118
rect 35420 16882 35476 17052
rect 35532 16996 35588 17006
rect 35532 16902 35588 16940
rect 35420 16830 35422 16882
rect 35474 16830 35476 16882
rect 35420 16818 35476 16830
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34860 16210 34916 16222
rect 34860 16158 34862 16210
rect 34914 16158 34916 16210
rect 34860 15876 34916 16158
rect 35532 16212 35588 16222
rect 35532 16118 35588 16156
rect 34860 15810 34916 15820
rect 34188 15092 34356 15148
rect 35644 15148 35700 27132
rect 36316 27076 36372 27086
rect 36316 26982 36372 27020
rect 35868 26962 35924 26974
rect 35868 26910 35870 26962
rect 35922 26910 35924 26962
rect 35756 26850 35812 26862
rect 35756 26798 35758 26850
rect 35810 26798 35812 26850
rect 35756 26516 35812 26798
rect 35868 26740 35924 26910
rect 35868 26674 35924 26684
rect 36204 26852 36260 26862
rect 35756 26460 36148 26516
rect 36092 26292 36148 26460
rect 36204 26514 36260 26796
rect 36204 26462 36206 26514
rect 36258 26462 36260 26514
rect 36204 26450 36260 26462
rect 36428 26516 36484 29932
rect 37100 29988 37156 31500
rect 37212 30212 37268 31612
rect 37436 31556 37492 32508
rect 38220 32452 38276 32462
rect 38220 32358 38276 32396
rect 37436 31490 37492 31500
rect 37996 31220 38052 31230
rect 37996 31126 38052 31164
rect 37548 30882 37604 30894
rect 37548 30830 37550 30882
rect 37602 30830 37604 30882
rect 37548 30436 37604 30830
rect 37548 30370 37604 30380
rect 37212 30146 37268 30156
rect 36652 27970 36708 27982
rect 36652 27918 36654 27970
rect 36706 27918 36708 27970
rect 36652 26908 36708 27918
rect 37100 27746 37156 29932
rect 38556 29988 38612 29998
rect 38556 29894 38612 29932
rect 37100 27694 37102 27746
rect 37154 27694 37156 27746
rect 36652 26852 36820 26908
rect 36428 26450 36484 26460
rect 36764 26402 36820 26852
rect 36764 26350 36766 26402
rect 36818 26350 36820 26402
rect 36540 26292 36596 26302
rect 36092 26290 36596 26292
rect 36092 26238 36542 26290
rect 36594 26238 36596 26290
rect 36092 26236 36596 26238
rect 36540 26226 36596 26236
rect 35756 25620 35812 25630
rect 35756 25526 35812 25564
rect 36316 25396 36372 25406
rect 36316 24834 36372 25340
rect 36316 24782 36318 24834
rect 36370 24782 36372 24834
rect 36316 24770 36372 24782
rect 36428 24724 36484 24734
rect 36428 24050 36484 24668
rect 36652 24724 36708 24734
rect 36764 24724 36820 26350
rect 37100 26852 37156 27694
rect 38668 27188 38724 35756
rect 39004 35812 39060 37772
rect 39004 35746 39060 35756
rect 38892 33460 38948 33470
rect 38892 33366 38948 33404
rect 38892 30210 38948 30222
rect 38892 30158 38894 30210
rect 38946 30158 38948 30210
rect 38892 29988 38948 30158
rect 38892 29922 38948 29932
rect 38780 28756 38836 28766
rect 38780 28084 38836 28700
rect 38780 28082 39172 28084
rect 38780 28030 38782 28082
rect 38834 28030 39172 28082
rect 38780 28028 39172 28030
rect 38780 28018 38836 28028
rect 39116 27970 39172 28028
rect 39116 27918 39118 27970
rect 39170 27918 39172 27970
rect 39116 27906 39172 27918
rect 37100 26292 37156 26796
rect 38444 27132 38724 27188
rect 37212 26292 37268 26302
rect 37100 26290 37268 26292
rect 37100 26238 37214 26290
rect 37266 26238 37268 26290
rect 37100 26236 37268 26238
rect 38444 26292 38500 27132
rect 39004 27074 39060 27086
rect 39004 27022 39006 27074
rect 39058 27022 39060 27074
rect 38556 26852 38612 26862
rect 38668 26852 38724 26862
rect 39004 26852 39060 27022
rect 38612 26850 39060 26852
rect 38612 26798 38670 26850
rect 38722 26798 39060 26850
rect 38612 26796 39060 26798
rect 38556 26786 38612 26796
rect 38668 26786 38724 26796
rect 38444 26236 38724 26292
rect 37212 26226 37268 26236
rect 36876 26180 36932 26190
rect 36876 26086 36932 26124
rect 37996 26180 38052 26190
rect 37996 26086 38052 26124
rect 36876 24724 36932 24734
rect 36652 24722 36876 24724
rect 36652 24670 36654 24722
rect 36706 24670 36876 24722
rect 36652 24668 36876 24670
rect 36652 24658 36708 24668
rect 36876 24658 36932 24668
rect 36652 24500 36708 24510
rect 36652 24406 36708 24444
rect 37772 24500 37828 24510
rect 36428 23998 36430 24050
rect 36482 23998 36484 24050
rect 36428 23940 36484 23998
rect 37772 24050 37828 24444
rect 37772 23998 37774 24050
rect 37826 23998 37828 24050
rect 37772 23986 37828 23998
rect 36428 23874 36484 23884
rect 37100 23940 37156 23950
rect 37100 23846 37156 23884
rect 37884 23940 37940 23950
rect 37884 21810 37940 23884
rect 37884 21758 37886 21810
rect 37938 21758 37940 21810
rect 37100 21084 37380 21140
rect 36988 20690 37044 20702
rect 36988 20638 36990 20690
rect 37042 20638 37044 20690
rect 35756 20580 35812 20590
rect 35756 20486 35812 20524
rect 36652 20580 36708 20590
rect 36988 20580 37044 20638
rect 36708 20524 37044 20580
rect 35756 20244 35812 20254
rect 35756 20130 35812 20188
rect 35756 20078 35758 20130
rect 35810 20078 35812 20130
rect 35756 20066 35812 20078
rect 36316 20018 36372 20030
rect 36316 19966 36318 20018
rect 36370 19966 36372 20018
rect 36316 19458 36372 19966
rect 36540 20020 36596 20030
rect 36540 19926 36596 19964
rect 36652 20020 36708 20524
rect 36764 20020 36820 20030
rect 36652 20018 36820 20020
rect 36652 19966 36766 20018
rect 36818 19966 36820 20018
rect 36652 19964 36820 19966
rect 36428 19908 36484 19918
rect 36428 19814 36484 19852
rect 36316 19406 36318 19458
rect 36370 19406 36372 19458
rect 36316 19394 36372 19406
rect 35980 19236 36036 19246
rect 35868 19012 35924 19022
rect 35868 18452 35924 18956
rect 35868 18386 35924 18396
rect 35980 17666 36036 19180
rect 36428 19236 36484 19246
rect 36428 19142 36484 19180
rect 36316 19012 36372 19022
rect 36316 18918 36372 18956
rect 35980 17614 35982 17666
rect 36034 17614 36036 17666
rect 35868 17444 35924 17454
rect 35756 16770 35812 16782
rect 35756 16718 35758 16770
rect 35810 16718 35812 16770
rect 35756 15428 35812 16718
rect 35756 15362 35812 15372
rect 35868 15316 35924 17388
rect 35980 17220 36036 17614
rect 36092 17444 36148 17454
rect 36092 17350 36148 17388
rect 36316 17442 36372 17454
rect 36316 17390 36318 17442
rect 36370 17390 36372 17442
rect 35980 17164 36148 17220
rect 35980 16882 36036 16894
rect 35980 16830 35982 16882
rect 36034 16830 36036 16882
rect 35980 16322 36036 16830
rect 35980 16270 35982 16322
rect 36034 16270 36036 16322
rect 35980 16258 36036 16270
rect 36092 16098 36148 17164
rect 36204 16996 36260 17006
rect 36316 16996 36372 17390
rect 36428 17108 36484 17118
rect 36652 17108 36708 19964
rect 36764 19954 36820 19964
rect 37100 19458 37156 21084
rect 37324 21028 37380 21084
rect 37324 20972 37604 21028
rect 37212 20916 37268 20926
rect 37268 20860 37380 20916
rect 37212 20850 37268 20860
rect 37212 20690 37268 20702
rect 37212 20638 37214 20690
rect 37266 20638 37268 20690
rect 37212 20244 37268 20638
rect 37212 20178 37268 20188
rect 37324 20020 37380 20860
rect 37548 20802 37604 20972
rect 37884 20916 37940 21758
rect 37940 20860 38276 20916
rect 37884 20850 37940 20860
rect 37548 20750 37550 20802
rect 37602 20750 37604 20802
rect 37548 20738 37604 20750
rect 38220 20802 38276 20860
rect 38220 20750 38222 20802
rect 38274 20750 38276 20802
rect 38220 20738 38276 20750
rect 37436 20692 37492 20702
rect 37436 20598 37492 20636
rect 37884 20356 37940 20366
rect 37324 20018 37716 20020
rect 37324 19966 37326 20018
rect 37378 19966 37716 20018
rect 37324 19964 37716 19966
rect 37324 19954 37380 19964
rect 37100 19406 37102 19458
rect 37154 19406 37156 19458
rect 37100 19394 37156 19406
rect 37212 19348 37268 19358
rect 36988 19236 37044 19246
rect 36988 19142 37044 19180
rect 37100 19124 37156 19134
rect 37212 19124 37268 19292
rect 37100 19122 37268 19124
rect 37100 19070 37102 19122
rect 37154 19070 37268 19122
rect 37100 19068 37268 19070
rect 37660 19346 37716 19964
rect 37660 19294 37662 19346
rect 37714 19294 37716 19346
rect 37100 19058 37156 19068
rect 37660 18562 37716 19294
rect 37660 18510 37662 18562
rect 37714 18510 37716 18562
rect 37100 17444 37156 17454
rect 37100 17350 37156 17388
rect 36484 17052 36708 17108
rect 36428 17042 36484 17052
rect 36204 16994 36372 16996
rect 36204 16942 36206 16994
rect 36258 16942 36372 16994
rect 36204 16940 36372 16942
rect 36204 16930 36260 16940
rect 36428 16884 36484 16894
rect 36428 16790 36484 16828
rect 36652 16882 36708 17052
rect 37660 17106 37716 18510
rect 37660 17054 37662 17106
rect 37714 17054 37716 17106
rect 36652 16830 36654 16882
rect 36706 16830 36708 16882
rect 36652 16818 36708 16830
rect 37212 16882 37268 16894
rect 37212 16830 37214 16882
rect 37266 16830 37268 16882
rect 36316 16772 36372 16782
rect 36316 16678 36372 16716
rect 37100 16324 37156 16334
rect 36092 16046 36094 16098
rect 36146 16046 36148 16098
rect 36092 16034 36148 16046
rect 36316 16212 36372 16222
rect 35868 15250 35924 15260
rect 35980 15876 36036 15886
rect 35644 15092 35924 15148
rect 34188 13076 34244 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35868 14308 35924 15092
rect 35868 14242 35924 14252
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34188 13010 34244 13020
rect 34860 13076 34916 13086
rect 34860 12982 34916 13020
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 33964 11506 34020 11676
rect 33964 11454 33966 11506
rect 34018 11454 34020 11506
rect 33964 11442 34020 11454
rect 34524 11172 34580 11182
rect 34524 11078 34580 11116
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35980 8932 36036 15820
rect 36316 15314 36372 16156
rect 36988 16212 37044 16222
rect 36988 16098 37044 16156
rect 36988 16046 36990 16098
rect 37042 16046 37044 16098
rect 36988 16034 37044 16046
rect 37100 15652 37156 16268
rect 37212 15876 37268 16830
rect 37660 16212 37716 17054
rect 37660 16146 37716 16156
rect 37772 16772 37828 16782
rect 37772 16210 37828 16716
rect 37772 16158 37774 16210
rect 37826 16158 37828 16210
rect 37772 16146 37828 16158
rect 37212 15810 37268 15820
rect 37100 15596 37268 15652
rect 37100 15428 37156 15438
rect 37100 15334 37156 15372
rect 36316 15262 36318 15314
rect 36370 15262 36372 15314
rect 36316 15250 36372 15262
rect 35980 8866 36036 8876
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35980 5012 36036 5022
rect 34188 4116 34244 4126
rect 34188 4022 34244 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 33628 3490 33684 3500
rect 33740 3444 33796 3454
rect 35532 3444 35588 3454
rect 33740 3350 33796 3388
rect 35196 3388 35532 3444
rect 35196 3332 35252 3388
rect 35532 3350 35588 3388
rect 35980 3442 36036 4956
rect 35980 3390 35982 3442
rect 36034 3390 36036 3442
rect 35980 3378 36036 3390
rect 36204 3554 36260 3566
rect 36204 3502 36206 3554
rect 36258 3502 36260 3554
rect 36204 3444 36260 3502
rect 36204 3378 36260 3388
rect 36988 3442 37044 3454
rect 36988 3390 36990 3442
rect 37042 3390 37044 3442
rect 34972 3276 35252 3332
rect 34972 800 35028 3276
rect 36988 3220 37044 3390
rect 37212 3442 37268 15596
rect 37884 15148 37940 20300
rect 37996 19908 38052 19918
rect 37996 19814 38052 19852
rect 38108 19348 38164 19358
rect 38108 19254 38164 19292
rect 38668 15876 38724 26236
rect 38892 25508 38948 25518
rect 38892 25414 38948 25452
rect 39116 25282 39172 25294
rect 39116 25230 39118 25282
rect 39170 25230 39172 25282
rect 39116 24834 39172 25230
rect 39116 24782 39118 24834
rect 39170 24782 39172 24834
rect 39116 24770 39172 24782
rect 39004 20692 39060 20702
rect 39004 20598 39060 20636
rect 39116 20244 39172 20254
rect 39116 17444 39172 20188
rect 39228 19908 39284 42476
rect 40236 42532 40292 42542
rect 40236 42438 40292 42476
rect 39788 41524 39844 41534
rect 39564 39620 39620 39630
rect 39564 39618 39732 39620
rect 39564 39566 39566 39618
rect 39618 39566 39732 39618
rect 39564 39564 39732 39566
rect 39564 39554 39620 39564
rect 39676 38612 39732 39564
rect 39788 39394 39844 41468
rect 39788 39342 39790 39394
rect 39842 39342 39844 39394
rect 39788 39330 39844 39342
rect 39676 38556 40180 38612
rect 40124 38274 40180 38556
rect 40124 38222 40126 38274
rect 40178 38222 40180 38274
rect 40124 38210 40180 38222
rect 39788 38052 39844 38062
rect 39788 37958 39844 37996
rect 39340 37940 39396 37950
rect 39340 35586 39396 37884
rect 39340 35534 39342 35586
rect 39394 35534 39396 35586
rect 39340 35140 39396 35534
rect 39340 35074 39396 35084
rect 40460 34914 40516 34926
rect 40460 34862 40462 34914
rect 40514 34862 40516 34914
rect 40124 34692 40180 34702
rect 40460 34692 40516 34862
rect 40124 34690 40516 34692
rect 40124 34638 40126 34690
rect 40178 34638 40516 34690
rect 40124 34636 40516 34638
rect 40124 33236 40180 34636
rect 40572 34580 40628 42588
rect 40796 42550 40852 42588
rect 40908 42532 40964 42702
rect 40908 42466 40964 42476
rect 41020 41524 41076 45054
rect 43148 45106 43876 45108
rect 43148 45054 43822 45106
rect 43874 45054 43876 45106
rect 43148 45052 43876 45054
rect 41580 44436 41636 44446
rect 41580 42978 41636 44380
rect 41580 42926 41582 42978
rect 41634 42926 41636 42978
rect 41580 42914 41636 42926
rect 41916 44212 41972 44222
rect 41916 42978 41972 44156
rect 42812 44212 42868 44222
rect 42812 44118 42868 44156
rect 43148 44210 43204 45052
rect 43820 45042 43876 45052
rect 43820 44324 43876 44334
rect 43148 44158 43150 44210
rect 43202 44158 43204 44210
rect 43148 44146 43204 44158
rect 43484 44210 43540 44222
rect 43484 44158 43486 44210
rect 43538 44158 43540 44210
rect 41916 42926 41918 42978
rect 41970 42926 41972 42978
rect 41916 42914 41972 42926
rect 41020 41458 41076 41468
rect 40684 37940 40740 37950
rect 40684 37846 40740 37884
rect 41132 37828 41188 37838
rect 41132 37734 41188 37772
rect 41020 36484 41076 36494
rect 41020 36482 41636 36484
rect 41020 36430 41022 36482
rect 41074 36430 41636 36482
rect 41020 36428 41636 36430
rect 41020 36418 41076 36428
rect 41244 36260 41300 36270
rect 41244 36166 41300 36204
rect 41244 36036 41300 36046
rect 41244 35138 41300 35980
rect 41244 35086 41246 35138
rect 41298 35086 41300 35138
rect 41244 35074 41300 35086
rect 41580 35138 41636 36428
rect 41580 35086 41582 35138
rect 41634 35086 41636 35138
rect 41580 35074 41636 35086
rect 40684 34804 40740 34814
rect 40684 34710 40740 34748
rect 41020 34804 41076 34814
rect 39676 30100 39732 30110
rect 39676 30006 39732 30044
rect 39564 28756 39620 28766
rect 39620 28700 39956 28756
rect 39564 28662 39620 28700
rect 39340 27970 39396 27982
rect 39340 27918 39342 27970
rect 39394 27918 39396 27970
rect 39340 26404 39396 27918
rect 39900 27970 39956 28700
rect 39900 27918 39902 27970
rect 39954 27918 39956 27970
rect 39900 27906 39956 27918
rect 40012 27746 40068 27758
rect 40012 27694 40014 27746
rect 40066 27694 40068 27746
rect 39452 27636 39508 27646
rect 39452 27634 39844 27636
rect 39452 27582 39454 27634
rect 39506 27582 39844 27634
rect 39452 27580 39844 27582
rect 39452 27570 39508 27580
rect 39788 27186 39844 27580
rect 39788 27134 39790 27186
rect 39842 27134 39844 27186
rect 39788 27122 39844 27134
rect 40012 26516 40068 27694
rect 39564 26460 40068 26516
rect 39340 26348 39508 26404
rect 39340 26068 39396 26078
rect 39340 25508 39396 26012
rect 39340 25414 39396 25452
rect 39452 25284 39508 26348
rect 39564 25506 39620 26460
rect 40124 25844 40180 33180
rect 40348 34524 40628 34580
rect 40348 32788 40404 34524
rect 40348 32450 40404 32732
rect 40348 32398 40350 32450
rect 40402 32398 40404 32450
rect 40348 32386 40404 32398
rect 41020 33458 41076 34748
rect 42140 34804 42196 34814
rect 42140 34710 42196 34748
rect 41020 33406 41022 33458
rect 41074 33406 41076 33458
rect 41020 32340 41076 33406
rect 41020 32274 41076 32284
rect 41132 31332 41188 31342
rect 40236 27860 40292 27898
rect 40236 27794 40292 27804
rect 39564 25454 39566 25506
rect 39618 25454 39620 25506
rect 39564 25442 39620 25454
rect 39900 25788 40180 25844
rect 40236 26964 40292 26974
rect 40236 26178 40292 26908
rect 40236 26126 40238 26178
rect 40290 26126 40292 26178
rect 39452 25228 39620 25284
rect 39340 24836 39396 24846
rect 39564 24836 39620 25228
rect 39676 24836 39732 24846
rect 39340 24834 39508 24836
rect 39340 24782 39342 24834
rect 39394 24782 39508 24834
rect 39340 24780 39508 24782
rect 39564 24834 39732 24836
rect 39564 24782 39678 24834
rect 39730 24782 39732 24834
rect 39564 24780 39732 24782
rect 39340 24770 39396 24780
rect 39452 24722 39508 24780
rect 39452 24670 39454 24722
rect 39506 24670 39508 24722
rect 39452 24658 39508 24670
rect 39676 24724 39732 24780
rect 39676 24658 39732 24668
rect 39788 24500 39844 24510
rect 39788 24406 39844 24444
rect 39900 24276 39956 25788
rect 39676 24220 39956 24276
rect 40012 25620 40068 25630
rect 39676 20244 39732 24220
rect 39900 24052 39956 24062
rect 40012 24052 40068 25564
rect 40124 25508 40180 25518
rect 40124 25414 40180 25452
rect 39900 24050 40068 24052
rect 39900 23998 39902 24050
rect 39954 23998 40068 24050
rect 39900 23996 40068 23998
rect 39900 20188 39956 23996
rect 40124 23940 40180 23950
rect 40124 23378 40180 23884
rect 40124 23326 40126 23378
rect 40178 23326 40180 23378
rect 40124 23314 40180 23326
rect 39676 20178 39732 20188
rect 39228 19012 39284 19852
rect 39228 18946 39284 18956
rect 39788 20132 39956 20188
rect 39116 17378 39172 17388
rect 38668 15810 38724 15820
rect 39228 15876 39284 15886
rect 37548 15092 37940 15148
rect 39228 15202 39284 15820
rect 39228 15150 39230 15202
rect 39282 15150 39284 15202
rect 39228 15138 39284 15150
rect 37548 8428 37604 15092
rect 37436 8372 37604 8428
rect 37436 5012 37492 8372
rect 37436 4946 37492 4956
rect 39788 5012 39844 20132
rect 40124 19908 40180 19918
rect 40124 19814 40180 19852
rect 39900 17444 39956 17454
rect 39956 17388 40068 17444
rect 39900 17378 39956 17388
rect 40012 16210 40068 17388
rect 40012 16158 40014 16210
rect 40066 16158 40068 16210
rect 40012 16146 40068 16158
rect 39900 16100 39956 16110
rect 39900 15538 39956 16044
rect 39900 15486 39902 15538
rect 39954 15486 39956 15538
rect 39900 15474 39956 15486
rect 39788 4946 39844 4956
rect 40236 4564 40292 26126
rect 40460 23940 40516 23950
rect 40460 23846 40516 23884
rect 41132 20914 41188 31276
rect 41692 31332 41748 31342
rect 41244 31220 41300 31230
rect 41244 31126 41300 31164
rect 41692 31218 41748 31276
rect 42364 31332 42420 31342
rect 41692 31166 41694 31218
rect 41746 31166 41748 31218
rect 41692 31154 41748 31166
rect 41804 31220 41860 31230
rect 41804 30322 41860 31164
rect 42364 30994 42420 31276
rect 42588 31220 42644 31230
rect 42588 31106 42644 31164
rect 43484 31218 43540 44158
rect 43820 44210 43876 44268
rect 43820 44158 43822 44210
rect 43874 44158 43876 44210
rect 43820 44146 43876 44158
rect 43932 36260 43988 45838
rect 44380 44548 44436 49200
rect 44604 46116 44660 46126
rect 44604 46022 44660 46060
rect 44828 45332 44884 45342
rect 44828 45238 44884 45276
rect 44380 44482 44436 44492
rect 44828 44324 44884 44334
rect 44828 44230 44884 44268
rect 45276 43650 45332 43662
rect 45276 43598 45278 43650
rect 45330 43598 45332 43650
rect 44940 43538 44996 43550
rect 44940 43486 44942 43538
rect 44994 43486 44996 43538
rect 44604 43428 44660 43438
rect 44940 43428 44996 43486
rect 44604 43426 44996 43428
rect 44604 43374 44606 43426
rect 44658 43374 44996 43426
rect 44604 43372 44996 43374
rect 44604 42868 44660 43372
rect 44604 42802 44660 42812
rect 45276 42756 45332 43598
rect 45612 43540 45668 43550
rect 45612 43446 45668 43484
rect 45724 43428 45780 49200
rect 45836 44548 45892 44558
rect 45836 44454 45892 44492
rect 45724 43362 45780 43372
rect 46620 43428 46676 43438
rect 46620 43334 46676 43372
rect 47068 42978 47124 49200
rect 48188 46452 48244 46462
rect 47628 46004 47684 46014
rect 48188 46004 48244 46396
rect 47628 46002 48244 46004
rect 47628 45950 47630 46002
rect 47682 45950 48244 46002
rect 47628 45948 48244 45950
rect 47628 45938 47684 45948
rect 48188 45890 48244 45948
rect 48188 45838 48190 45890
rect 48242 45838 48244 45890
rect 48188 45826 48244 45838
rect 47852 45666 47908 45678
rect 47852 45614 47854 45666
rect 47906 45614 47908 45666
rect 47852 44436 47908 45614
rect 47852 44370 47908 44380
rect 47068 42926 47070 42978
rect 47122 42926 47124 42978
rect 47068 42914 47124 42926
rect 45612 42756 45668 42766
rect 45276 42754 45668 42756
rect 45276 42702 45614 42754
rect 45666 42702 45668 42754
rect 45276 42700 45668 42702
rect 45612 42690 45668 42700
rect 47628 41076 47684 41086
rect 47628 40982 47684 41020
rect 48188 41076 48244 41086
rect 48188 40982 48244 41020
rect 47852 40962 47908 40974
rect 47852 40910 47854 40962
rect 47906 40910 47908 40962
rect 46172 38724 46228 38734
rect 43932 36194 43988 36204
rect 44492 37268 44548 37278
rect 43484 31166 43486 31218
rect 43538 31166 43540 31218
rect 43484 31154 43540 31166
rect 42588 31054 42590 31106
rect 42642 31054 42644 31106
rect 42588 31042 42644 31054
rect 43148 31108 43204 31118
rect 42364 30942 42366 30994
rect 42418 30942 42420 30994
rect 42364 30930 42420 30942
rect 43148 30994 43204 31052
rect 43148 30942 43150 30994
rect 43202 30942 43204 30994
rect 43148 30930 43204 30942
rect 41804 30270 41806 30322
rect 41858 30270 41860 30322
rect 41804 30258 41860 30270
rect 42028 30324 42084 30334
rect 41916 27860 41972 27870
rect 41916 27186 41972 27804
rect 41916 27134 41918 27186
rect 41970 27134 41972 27186
rect 41916 27122 41972 27134
rect 42028 25508 42084 30268
rect 42028 25442 42084 25452
rect 43372 25396 43428 25406
rect 41244 24500 41300 24510
rect 41244 24050 41300 24444
rect 41244 23998 41246 24050
rect 41298 23998 41300 24050
rect 41244 23986 41300 23998
rect 43372 24050 43428 25340
rect 43372 23998 43374 24050
rect 43426 23998 43428 24050
rect 41132 20862 41134 20914
rect 41186 20862 41188 20914
rect 41132 19348 41188 20862
rect 43372 20188 43428 23998
rect 43372 20132 43540 20188
rect 41132 19282 41188 19292
rect 42028 5012 42084 5022
rect 40348 4564 40404 4574
rect 40236 4508 40348 4564
rect 40348 4470 40404 4508
rect 41244 4564 41300 4574
rect 41244 4338 41300 4508
rect 41244 4286 41246 4338
rect 41298 4286 41300 4338
rect 41244 4274 41300 4286
rect 41020 4116 41076 4126
rect 39004 3668 39060 3678
rect 37212 3390 37214 3442
rect 37266 3390 37268 3442
rect 37212 3378 37268 3390
rect 37436 3554 37492 3566
rect 37436 3502 37438 3554
rect 37490 3502 37492 3554
rect 37436 3220 37492 3502
rect 36988 3164 37492 3220
rect 36988 800 37044 3164
rect 39004 800 39060 3612
rect 40012 3668 40068 3678
rect 40012 3574 40068 3612
rect 41020 800 41076 4060
rect 42028 3668 42084 4956
rect 42252 4116 42308 4126
rect 42252 4022 42308 4060
rect 42028 3554 42084 3612
rect 42812 3668 42868 3678
rect 42812 3574 42868 3612
rect 42028 3502 42030 3554
rect 42082 3502 42084 3554
rect 42028 3490 42084 3502
rect 43484 3556 43540 20132
rect 44492 4564 44548 37212
rect 44492 4498 44548 4508
rect 45052 25284 45108 25294
rect 43820 3668 43876 3678
rect 43484 3490 43540 3500
rect 43596 3666 43876 3668
rect 43596 3614 43822 3666
rect 43874 3614 43876 3666
rect 43596 3612 43876 3614
rect 43596 980 43652 3612
rect 43820 3602 43876 3612
rect 43036 924 43652 980
rect 43036 800 43092 924
rect 45052 800 45108 25228
rect 46172 20132 46228 38668
rect 47852 38052 47908 40910
rect 47852 37986 47908 37996
rect 47628 36372 47684 36382
rect 47628 36278 47684 36316
rect 48188 36372 48244 36382
rect 47852 36260 47908 36270
rect 47852 36166 47908 36204
rect 48188 35700 48244 36316
rect 48188 35634 48244 35644
rect 47852 31108 47908 31118
rect 47852 31014 47908 31052
rect 48188 30994 48244 31006
rect 48188 30942 48190 30994
rect 48242 30942 48244 30994
rect 47628 30884 47684 30894
rect 48188 30884 48244 30942
rect 47628 30882 48244 30884
rect 47628 30830 47630 30882
rect 47682 30830 48244 30882
rect 47628 30828 48244 30830
rect 47628 30818 47684 30828
rect 48188 30324 48244 30828
rect 48188 30258 48244 30268
rect 47852 25508 47908 25518
rect 47852 25394 47908 25452
rect 47852 25342 47854 25394
rect 47906 25342 47908 25394
rect 47852 25330 47908 25342
rect 48188 25394 48244 25406
rect 48188 25342 48190 25394
rect 48242 25342 48244 25394
rect 47628 25284 47684 25294
rect 47628 25190 47684 25228
rect 48188 25284 48244 25342
rect 48188 24948 48244 25228
rect 48188 24882 48244 24892
rect 46172 20066 46228 20076
rect 46284 21588 46340 21598
rect 46284 3668 46340 21532
rect 47852 20132 47908 20142
rect 47852 20038 47908 20076
rect 48188 20018 48244 20030
rect 48188 19966 48190 20018
rect 48242 19966 48244 20018
rect 47628 19908 47684 19918
rect 48188 19908 48244 19966
rect 47628 19906 48244 19908
rect 47628 19854 47630 19906
rect 47682 19854 48244 19906
rect 47628 19852 48244 19854
rect 47628 19842 47684 19852
rect 48188 19572 48244 19852
rect 48188 19506 48244 19516
rect 48188 14418 48244 14430
rect 48188 14366 48190 14418
rect 48242 14366 48244 14418
rect 47628 14306 47684 14318
rect 47628 14254 47630 14306
rect 47682 14254 47684 14306
rect 47628 14196 47684 14254
rect 47852 14308 47908 14318
rect 47852 14214 47908 14252
rect 47628 14130 47684 14140
rect 48188 14196 48244 14366
rect 48188 14130 48244 14140
rect 47852 9156 47908 9166
rect 47852 9062 47908 9100
rect 48188 9042 48244 9054
rect 48188 8990 48190 9042
rect 48242 8990 48244 9042
rect 47628 8930 47684 8942
rect 47628 8878 47630 8930
rect 47682 8878 47684 8930
rect 47628 8820 47684 8878
rect 47628 8754 47684 8764
rect 48188 8820 48244 8990
rect 48188 8754 48244 8764
rect 47852 4564 47908 4574
rect 47852 4470 47908 4508
rect 48188 4338 48244 4350
rect 48188 4286 48190 4338
rect 48242 4286 48244 4338
rect 46956 4228 47012 4238
rect 47628 4228 47684 4238
rect 48188 4228 48244 4286
rect 46956 4226 47124 4228
rect 46956 4174 46958 4226
rect 47010 4174 47124 4226
rect 46956 4172 47124 4174
rect 46956 4162 47012 4172
rect 46284 3602 46340 3612
rect 45724 3556 45780 3566
rect 45724 3462 45780 3500
rect 46620 3556 46676 3566
rect 46620 3462 46676 3500
rect 47068 2548 47124 4172
rect 47628 4226 48244 4228
rect 47628 4174 47630 4226
rect 47682 4174 48244 4226
rect 47628 4172 48244 4174
rect 47628 4162 47684 4172
rect 47852 3668 47908 3678
rect 47852 3574 47908 3612
rect 47404 3442 47460 3454
rect 47404 3390 47406 3442
rect 47458 3390 47460 3442
rect 47404 2548 47460 3390
rect 48188 3444 48244 4172
rect 48188 3378 48244 3388
rect 47068 2492 47460 2548
rect 47068 800 47124 2492
rect 2688 0 2800 800
rect 4704 0 4816 800
rect 6720 0 6832 800
rect 8736 0 8848 800
rect 10752 0 10864 800
rect 12768 0 12880 800
rect 14784 0 14896 800
rect 16800 0 16912 800
rect 18816 0 18928 800
rect 20832 0 20944 800
rect 22848 0 22960 800
rect 24864 0 24976 800
rect 26880 0 26992 800
rect 28896 0 29008 800
rect 30912 0 31024 800
rect 32928 0 33040 800
rect 34944 0 35056 800
rect 36960 0 37072 800
rect 38976 0 39088 800
rect 40992 0 41104 800
rect 43008 0 43120 800
rect 45024 0 45136 800
rect 47040 0 47152 800
<< via2 >>
rect 2716 46844 2772 46900
rect 1932 46002 1988 46004
rect 1932 45950 1934 46002
rect 1934 45950 1986 46002
rect 1986 45950 1988 46002
rect 1932 45948 1988 45950
rect 1820 44380 1876 44436
rect 1596 44268 1652 44324
rect 1484 43820 1540 43876
rect 1484 29820 1540 29876
rect 1932 42812 1988 42868
rect 2044 41356 2100 41412
rect 2156 42812 2212 42868
rect 2044 40908 2100 40964
rect 1932 39676 1988 39732
rect 1932 38108 1988 38164
rect 4844 47516 4900 47572
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4732 45890 4788 45892
rect 4732 45838 4734 45890
rect 4734 45838 4786 45890
rect 4786 45838 4788 45890
rect 4732 45836 4788 45838
rect 4284 45500 4340 45556
rect 5404 45836 5460 45892
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 3948 42588 4004 42644
rect 3836 40908 3892 40964
rect 2156 38108 2212 38164
rect 2828 38162 2884 38164
rect 2828 38110 2830 38162
rect 2830 38110 2882 38162
rect 2882 38110 2884 38162
rect 2828 38108 2884 38110
rect 3836 38668 3892 38724
rect 3276 38050 3332 38052
rect 3276 37998 3278 38050
rect 3278 37998 3330 38050
rect 3330 37998 3332 38050
rect 3276 37996 3332 37998
rect 2380 37266 2436 37268
rect 2380 37214 2382 37266
rect 2382 37214 2434 37266
rect 2434 37214 2436 37266
rect 2380 37212 2436 37214
rect 2940 36652 2996 36708
rect 1932 36594 1988 36596
rect 1932 36542 1934 36594
rect 1934 36542 1986 36594
rect 1986 36542 1988 36594
rect 1932 36540 1988 36542
rect 3052 35868 3108 35924
rect 1932 34972 1988 35028
rect 2044 35420 2100 35476
rect 3612 37548 3668 37604
rect 3500 35868 3556 35924
rect 3164 34972 3220 35028
rect 2828 34914 2884 34916
rect 2828 34862 2830 34914
rect 2830 34862 2882 34914
rect 2882 34862 2884 34914
rect 2828 34860 2884 34862
rect 2940 34802 2996 34804
rect 2940 34750 2942 34802
rect 2942 34750 2994 34802
rect 2994 34750 2996 34802
rect 2940 34748 2996 34750
rect 2716 34188 2772 34244
rect 3052 34188 3108 34244
rect 1708 33404 1764 33460
rect 2492 33404 2548 33460
rect 1820 31836 1876 31892
rect 1932 31724 1988 31780
rect 1932 30322 1988 30324
rect 1932 30270 1934 30322
rect 1934 30270 1986 30322
rect 1986 30270 1988 30322
rect 1932 30268 1988 30270
rect 1932 28700 1988 28756
rect 2156 28754 2212 28756
rect 2156 28702 2158 28754
rect 2158 28702 2210 28754
rect 2210 28702 2212 28754
rect 2156 28700 2212 28702
rect 2940 27580 2996 27636
rect 1596 26460 1652 26516
rect 1932 27132 1988 27188
rect 2156 26908 2212 26964
rect 1932 25618 1988 25620
rect 1932 25566 1934 25618
rect 1934 25566 1986 25618
rect 1986 25566 1988 25618
rect 1932 25564 1988 25566
rect 2828 24610 2884 24612
rect 2828 24558 2830 24610
rect 2830 24558 2882 24610
rect 2882 24558 2884 24610
rect 2828 24556 2884 24558
rect 1932 24050 1988 24052
rect 1932 23998 1934 24050
rect 1934 23998 1986 24050
rect 1986 23998 1988 24050
rect 1932 23996 1988 23998
rect 2044 23100 2100 23156
rect 1932 22428 1988 22484
rect 1932 20914 1988 20916
rect 1932 20862 1934 20914
rect 1934 20862 1986 20914
rect 1986 20862 1988 20914
rect 1932 20860 1988 20862
rect 2268 20748 2324 20804
rect 1708 19852 1764 19908
rect 2492 19906 2548 19908
rect 2492 19854 2494 19906
rect 2494 19854 2546 19906
rect 2546 19854 2548 19906
rect 2492 19852 2548 19854
rect 2044 19740 2100 19796
rect 1708 19292 1764 19348
rect 1932 19068 1988 19124
rect 1708 18284 1764 18340
rect 1708 17724 1764 17780
rect 1820 16210 1876 16212
rect 1820 16158 1822 16210
rect 1822 16158 1874 16210
rect 1874 16158 1876 16210
rect 1820 16156 1876 16158
rect 1708 14588 1764 14644
rect 1820 13074 1876 13076
rect 1820 13022 1822 13074
rect 1822 13022 1874 13074
rect 1874 13022 1876 13074
rect 1820 13020 1876 13022
rect 1820 11506 1876 11508
rect 1820 11454 1822 11506
rect 1822 11454 1874 11506
rect 1874 11454 1876 11506
rect 1820 11452 1876 11454
rect 1820 9938 1876 9940
rect 1820 9886 1822 9938
rect 1822 9886 1874 9938
rect 1874 9886 1876 9938
rect 1820 9884 1876 9886
rect 2716 18956 2772 19012
rect 2492 18338 2548 18340
rect 2492 18286 2494 18338
rect 2494 18286 2546 18338
rect 2546 18286 2548 18338
rect 2492 18284 2548 18286
rect 2044 18172 2100 18228
rect 2268 17388 2324 17444
rect 2492 16828 2548 16884
rect 2604 16268 2660 16324
rect 2268 14140 2324 14196
rect 2044 9266 2100 9268
rect 2044 9214 2046 9266
rect 2046 9214 2098 9266
rect 2098 9214 2100 9266
rect 2044 9212 2100 9214
rect 2268 13746 2324 13748
rect 2268 13694 2270 13746
rect 2270 13694 2322 13746
rect 2322 13694 2324 13746
rect 2268 13692 2324 13694
rect 2268 12066 2324 12068
rect 2268 12014 2270 12066
rect 2270 12014 2322 12066
rect 2322 12014 2324 12066
rect 2268 12012 2324 12014
rect 2380 11452 2436 11508
rect 2268 10722 2324 10724
rect 2268 10670 2270 10722
rect 2270 10670 2322 10722
rect 2322 10670 2324 10722
rect 2268 10668 2324 10670
rect 1708 8316 1764 8372
rect 1708 7308 1764 7364
rect 1708 6748 1764 6804
rect 2492 8316 2548 8372
rect 2492 7362 2548 7364
rect 2492 7310 2494 7362
rect 2494 7310 2546 7362
rect 2546 7310 2548 7362
rect 2492 7308 2548 7310
rect 1820 5234 1876 5236
rect 1820 5182 1822 5234
rect 1822 5182 1874 5234
rect 1874 5182 1876 5234
rect 1820 5180 1876 5182
rect 1708 4172 1764 4228
rect 1708 3612 1764 3668
rect 2940 17554 2996 17556
rect 2940 17502 2942 17554
rect 2942 17502 2994 17554
rect 2994 17502 2996 17554
rect 2940 17500 2996 17502
rect 3612 34914 3668 34916
rect 3612 34862 3614 34914
rect 3614 34862 3666 34914
rect 3666 34862 3668 34914
rect 3612 34860 3668 34862
rect 3164 23212 3220 23268
rect 3612 33964 3668 34020
rect 4284 44044 4340 44100
rect 4844 44322 4900 44324
rect 4844 44270 4846 44322
rect 4846 44270 4898 44322
rect 4898 44270 4900 44322
rect 4844 44268 4900 44270
rect 4956 43932 5012 43988
rect 5628 46844 5684 46900
rect 5628 45948 5684 46004
rect 6636 46002 6692 46004
rect 6636 45950 6638 46002
rect 6638 45950 6690 46002
rect 6690 45950 6692 46002
rect 6636 45948 6692 45950
rect 5628 44268 5684 44324
rect 5964 44322 6020 44324
rect 5964 44270 5966 44322
rect 5966 44270 6018 44322
rect 6018 44270 6020 44322
rect 5964 44268 6020 44270
rect 5628 43708 5684 43764
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4284 42754 4340 42756
rect 4284 42702 4286 42754
rect 4286 42702 4338 42754
rect 4338 42702 4340 42754
rect 4284 42700 4340 42702
rect 4508 41858 4564 41860
rect 4508 41806 4510 41858
rect 4510 41806 4562 41858
rect 4562 41806 4564 41858
rect 4508 41804 4564 41806
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4844 41298 4900 41300
rect 4844 41246 4846 41298
rect 4846 41246 4898 41298
rect 4898 41246 4900 41298
rect 4844 41244 4900 41246
rect 4284 40236 4340 40292
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4844 38722 4900 38724
rect 4844 38670 4846 38722
rect 4846 38670 4898 38722
rect 4898 38670 4900 38722
rect 4844 38668 4900 38670
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5516 41244 5572 41300
rect 5292 39452 5348 39508
rect 4956 38108 5012 38164
rect 4284 37996 4340 38052
rect 4060 36540 4116 36596
rect 4284 37100 4340 37156
rect 4508 36988 4564 37044
rect 4844 37938 4900 37940
rect 4844 37886 4846 37938
rect 4846 37886 4898 37938
rect 4898 37886 4900 37938
rect 4844 37884 4900 37886
rect 4844 37548 4900 37604
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4844 36764 4900 36820
rect 5180 37436 5236 37492
rect 5180 36988 5236 37044
rect 4956 36428 5012 36484
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4284 35084 4340 35140
rect 5068 36370 5124 36372
rect 5068 36318 5070 36370
rect 5070 36318 5122 36370
rect 5122 36318 5124 36370
rect 5068 36316 5124 36318
rect 5628 40908 5684 40964
rect 5628 37266 5684 37268
rect 5628 37214 5630 37266
rect 5630 37214 5682 37266
rect 5682 37214 5684 37266
rect 5628 37212 5684 37214
rect 5628 36764 5684 36820
rect 5852 36652 5908 36708
rect 5740 36594 5796 36596
rect 5740 36542 5742 36594
rect 5742 36542 5794 36594
rect 5794 36542 5796 36594
rect 5740 36540 5796 36542
rect 6076 36482 6132 36484
rect 6076 36430 6078 36482
rect 6078 36430 6130 36482
rect 6130 36430 6132 36482
rect 6076 36428 6132 36430
rect 5516 36316 5572 36372
rect 7196 45612 7252 45668
rect 8428 45666 8484 45668
rect 8428 45614 8430 45666
rect 8430 45614 8482 45666
rect 8482 45614 8484 45666
rect 8428 45612 8484 45614
rect 7868 45218 7924 45220
rect 7868 45166 7870 45218
rect 7870 45166 7922 45218
rect 7922 45166 7924 45218
rect 7868 45164 7924 45166
rect 8652 45218 8708 45220
rect 8652 45166 8654 45218
rect 8654 45166 8706 45218
rect 8706 45166 8708 45218
rect 8652 45164 8708 45166
rect 8092 44380 8148 44436
rect 7420 43932 7476 43988
rect 6748 42700 6804 42756
rect 6972 41244 7028 41300
rect 6860 40962 6916 40964
rect 6860 40910 6862 40962
rect 6862 40910 6914 40962
rect 6914 40910 6916 40962
rect 6860 40908 6916 40910
rect 6636 40460 6692 40516
rect 7084 40514 7140 40516
rect 7084 40462 7086 40514
rect 7086 40462 7138 40514
rect 7138 40462 7140 40514
rect 7084 40460 7140 40462
rect 7308 41970 7364 41972
rect 7308 41918 7310 41970
rect 7310 41918 7362 41970
rect 7362 41918 7364 41970
rect 7308 41916 7364 41918
rect 7420 41858 7476 41860
rect 7420 41806 7422 41858
rect 7422 41806 7474 41858
rect 7474 41806 7476 41858
rect 7420 41804 7476 41806
rect 6748 40236 6804 40292
rect 7196 39900 7252 39956
rect 7308 39618 7364 39620
rect 7308 39566 7310 39618
rect 7310 39566 7362 39618
rect 7362 39566 7364 39618
rect 7308 39564 7364 39566
rect 6748 39506 6804 39508
rect 6748 39454 6750 39506
rect 6750 39454 6802 39506
rect 6802 39454 6804 39506
rect 6748 39452 6804 39454
rect 6188 35756 6244 35812
rect 4396 34802 4452 34804
rect 4396 34750 4398 34802
rect 4398 34750 4450 34802
rect 4450 34750 4452 34802
rect 4396 34748 4452 34750
rect 6636 34972 6692 35028
rect 4844 34748 4900 34804
rect 5628 34802 5684 34804
rect 5628 34750 5630 34802
rect 5630 34750 5682 34802
rect 5682 34750 5684 34802
rect 5628 34748 5684 34750
rect 5964 34802 6020 34804
rect 5964 34750 5966 34802
rect 5966 34750 6018 34802
rect 6018 34750 6020 34802
rect 5964 34748 6020 34750
rect 4508 34018 4564 34020
rect 4508 33966 4510 34018
rect 4510 33966 4562 34018
rect 4562 33966 4564 34018
rect 4508 33964 4564 33966
rect 3388 16882 3444 16884
rect 3388 16830 3390 16882
rect 3390 16830 3442 16882
rect 3442 16830 3444 16882
rect 3388 16828 3444 16830
rect 4060 31666 4116 31668
rect 4060 31614 4062 31666
rect 4062 31614 4114 31666
rect 4114 31614 4116 31666
rect 4060 31612 4116 31614
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 6412 33740 6468 33796
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4284 31724 4340 31780
rect 5068 31836 5124 31892
rect 3948 30882 4004 30884
rect 3948 30830 3950 30882
rect 3950 30830 4002 30882
rect 4002 30830 4004 30882
rect 3948 30828 4004 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4172 28812 4228 28868
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4284 28700 4340 28756
rect 5740 31778 5796 31780
rect 5740 31726 5742 31778
rect 5742 31726 5794 31778
rect 5794 31726 5796 31778
rect 5740 31724 5796 31726
rect 5852 31554 5908 31556
rect 5852 31502 5854 31554
rect 5854 31502 5906 31554
rect 5906 31502 5908 31554
rect 5852 31500 5908 31502
rect 6076 31164 6132 31220
rect 4060 27804 4116 27860
rect 5068 28028 5124 28084
rect 4284 27580 4340 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4508 26908 4564 26964
rect 4956 26124 5012 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 7308 35308 7364 35364
rect 7308 35138 7364 35140
rect 7308 35086 7310 35138
rect 7310 35086 7362 35138
rect 7362 35086 7364 35138
rect 7308 35084 7364 35086
rect 7756 42642 7812 42644
rect 7756 42590 7758 42642
rect 7758 42590 7810 42642
rect 7810 42590 7812 42642
rect 7756 42588 7812 42590
rect 7644 42476 7700 42532
rect 8092 43932 8148 43988
rect 8092 42812 8148 42868
rect 8092 42642 8148 42644
rect 8092 42590 8094 42642
rect 8094 42590 8146 42642
rect 8146 42590 8148 42642
rect 8092 42588 8148 42590
rect 9324 43596 9380 43652
rect 8988 42812 9044 42868
rect 8764 42754 8820 42756
rect 8764 42702 8766 42754
rect 8766 42702 8818 42754
rect 8818 42702 8820 42754
rect 8764 42700 8820 42702
rect 8428 42530 8484 42532
rect 8428 42478 8430 42530
rect 8430 42478 8482 42530
rect 8482 42478 8484 42530
rect 8428 42476 8484 42478
rect 8092 42364 8148 42420
rect 8428 42082 8484 42084
rect 8428 42030 8430 42082
rect 8430 42030 8482 42082
rect 8482 42030 8484 42082
rect 8428 42028 8484 42030
rect 9436 43372 9492 43428
rect 8988 42476 9044 42532
rect 8652 41970 8708 41972
rect 8652 41918 8654 41970
rect 8654 41918 8706 41970
rect 8706 41918 8708 41970
rect 8652 41916 8708 41918
rect 8204 41804 8260 41860
rect 8204 39900 8260 39956
rect 9324 42028 9380 42084
rect 8876 41244 8932 41300
rect 9212 41298 9268 41300
rect 9212 41246 9214 41298
rect 9214 41246 9266 41298
rect 9266 41246 9268 41298
rect 9212 41244 9268 41246
rect 8988 41132 9044 41188
rect 8428 40684 8484 40740
rect 8988 40684 9044 40740
rect 8428 40348 8484 40404
rect 8988 40348 9044 40404
rect 8540 39004 8596 39060
rect 7644 37996 7700 38052
rect 7756 37100 7812 37156
rect 8092 37436 8148 37492
rect 8092 36988 8148 37044
rect 8316 36428 8372 36484
rect 7980 34748 8036 34804
rect 7420 33740 7476 33796
rect 7644 33964 7700 34020
rect 6636 31836 6692 31892
rect 6412 24892 6468 24948
rect 6524 30380 6580 30436
rect 4284 24556 4340 24612
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 5964 23548 6020 23604
rect 4284 23212 4340 23268
rect 5740 23266 5796 23268
rect 5740 23214 5742 23266
rect 5742 23214 5794 23266
rect 5794 23214 5796 23266
rect 5740 23212 5796 23214
rect 5852 23154 5908 23156
rect 5852 23102 5854 23154
rect 5854 23102 5906 23154
rect 5906 23102 5908 23154
rect 5852 23100 5908 23102
rect 5180 23042 5236 23044
rect 5180 22990 5182 23042
rect 5182 22990 5234 23042
rect 5234 22990 5236 23042
rect 5180 22988 5236 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4508 22540 4564 22596
rect 4172 22482 4228 22484
rect 4172 22430 4174 22482
rect 4174 22430 4226 22482
rect 4226 22430 4228 22482
rect 4172 22428 4228 22430
rect 6860 27298 6916 27300
rect 6860 27246 6862 27298
rect 6862 27246 6914 27298
rect 6914 27246 6916 27298
rect 6860 27244 6916 27246
rect 6748 26962 6804 26964
rect 6748 26910 6750 26962
rect 6750 26910 6802 26962
rect 6802 26910 6804 26962
rect 6748 26908 6804 26910
rect 7980 33292 8036 33348
rect 8428 36370 8484 36372
rect 8428 36318 8430 36370
rect 8430 36318 8482 36370
rect 8482 36318 8484 36370
rect 8428 36316 8484 36318
rect 8316 35308 8372 35364
rect 8876 37100 8932 37156
rect 8540 34972 8596 35028
rect 9548 42588 9604 42644
rect 9436 39004 9492 39060
rect 9660 42476 9716 42532
rect 8204 31948 8260 32004
rect 7644 31388 7700 31444
rect 7980 31612 8036 31668
rect 8092 31500 8148 31556
rect 8316 31554 8372 31556
rect 8316 31502 8318 31554
rect 8318 31502 8370 31554
rect 8370 31502 8372 31554
rect 8316 31500 8372 31502
rect 8540 31554 8596 31556
rect 8540 31502 8542 31554
rect 8542 31502 8594 31554
rect 8594 31502 8596 31554
rect 8540 31500 8596 31502
rect 9548 37378 9604 37380
rect 9548 37326 9550 37378
rect 9550 37326 9602 37378
rect 9602 37326 9604 37378
rect 9548 37324 9604 37326
rect 9548 37100 9604 37156
rect 10556 43650 10612 43652
rect 10556 43598 10558 43650
rect 10558 43598 10610 43650
rect 10610 43598 10612 43650
rect 10556 43596 10612 43598
rect 9884 42588 9940 42644
rect 9996 42700 10052 42756
rect 9996 42082 10052 42084
rect 9996 42030 9998 42082
rect 9998 42030 10050 42082
rect 10050 42030 10052 42082
rect 9996 42028 10052 42030
rect 11116 43036 11172 43092
rect 10668 41916 10724 41972
rect 10780 41356 10836 41412
rect 10892 41692 10948 41748
rect 10668 40460 10724 40516
rect 10220 39564 10276 39620
rect 9884 38834 9940 38836
rect 9884 38782 9886 38834
rect 9886 38782 9938 38834
rect 9938 38782 9940 38834
rect 9884 38780 9940 38782
rect 10556 38834 10612 38836
rect 10556 38782 10558 38834
rect 10558 38782 10610 38834
rect 10610 38782 10612 38834
rect 10556 38780 10612 38782
rect 9996 38220 10052 38276
rect 10444 38108 10500 38164
rect 9996 37324 10052 37380
rect 9772 37100 9828 37156
rect 9884 36428 9940 36484
rect 10220 37212 10276 37268
rect 9212 32284 9268 32340
rect 9884 35698 9940 35700
rect 9884 35646 9886 35698
rect 9886 35646 9938 35698
rect 9938 35646 9940 35698
rect 9884 35644 9940 35646
rect 9436 34802 9492 34804
rect 9436 34750 9438 34802
rect 9438 34750 9490 34802
rect 9490 34750 9492 34802
rect 9436 34748 9492 34750
rect 10892 39564 10948 39620
rect 10668 36876 10724 36932
rect 10332 35868 10388 35924
rect 10668 35644 10724 35700
rect 9660 35196 9716 35252
rect 9772 35084 9828 35140
rect 9548 33346 9604 33348
rect 9548 33294 9550 33346
rect 9550 33294 9602 33346
rect 9602 33294 9604 33346
rect 9548 33292 9604 33294
rect 9772 33292 9828 33348
rect 10108 33292 10164 33348
rect 9884 33068 9940 33124
rect 9436 31948 9492 32004
rect 8876 31500 8932 31556
rect 8764 31276 8820 31332
rect 9100 31052 9156 31108
rect 7756 30994 7812 30996
rect 7756 30942 7758 30994
rect 7758 30942 7810 30994
rect 7810 30942 7812 30994
rect 7756 30940 7812 30942
rect 7644 30882 7700 30884
rect 7644 30830 7646 30882
rect 7646 30830 7698 30882
rect 7698 30830 7700 30882
rect 7644 30828 7700 30830
rect 7980 30268 8036 30324
rect 7532 28754 7588 28756
rect 7532 28702 7534 28754
rect 7534 28702 7586 28754
rect 7586 28702 7588 28754
rect 7532 28700 7588 28702
rect 7644 28642 7700 28644
rect 7644 28590 7646 28642
rect 7646 28590 7698 28642
rect 7698 28590 7700 28642
rect 7644 28588 7700 28590
rect 7644 27804 7700 27860
rect 7756 27746 7812 27748
rect 7756 27694 7758 27746
rect 7758 27694 7810 27746
rect 7810 27694 7812 27746
rect 7756 27692 7812 27694
rect 7420 26796 7476 26852
rect 8540 30882 8596 30884
rect 8540 30830 8542 30882
rect 8542 30830 8594 30882
rect 8594 30830 8596 30882
rect 8540 30828 8596 30830
rect 8316 30268 8372 30324
rect 8764 30268 8820 30324
rect 9884 31948 9940 32004
rect 10108 31890 10164 31892
rect 10108 31838 10110 31890
rect 10110 31838 10162 31890
rect 10162 31838 10164 31890
rect 10108 31836 10164 31838
rect 9548 31724 9604 31780
rect 9324 31612 9380 31668
rect 9660 31666 9716 31668
rect 9660 31614 9662 31666
rect 9662 31614 9714 31666
rect 9714 31614 9716 31666
rect 9660 31612 9716 31614
rect 9772 31554 9828 31556
rect 9772 31502 9774 31554
rect 9774 31502 9826 31554
rect 9826 31502 9828 31554
rect 9772 31500 9828 31502
rect 11116 38162 11172 38164
rect 11116 38110 11118 38162
rect 11118 38110 11170 38162
rect 11170 38110 11172 38162
rect 11116 38108 11172 38110
rect 10892 37266 10948 37268
rect 10892 37214 10894 37266
rect 10894 37214 10946 37266
rect 10946 37214 10948 37266
rect 10892 37212 10948 37214
rect 11116 36594 11172 36596
rect 11116 36542 11118 36594
rect 11118 36542 11170 36594
rect 11170 36542 11172 36594
rect 11116 36540 11172 36542
rect 11676 45500 11732 45556
rect 11340 44268 11396 44324
rect 16380 45836 16436 45892
rect 17052 45890 17108 45892
rect 17052 45838 17054 45890
rect 17054 45838 17106 45890
rect 17106 45838 17108 45890
rect 17052 45836 17108 45838
rect 11340 43372 11396 43428
rect 12012 43596 12068 43652
rect 11564 42812 11620 42868
rect 12684 42866 12740 42868
rect 12684 42814 12686 42866
rect 12686 42814 12738 42866
rect 12738 42814 12740 42866
rect 12684 42812 12740 42814
rect 11452 42028 11508 42084
rect 11340 41692 11396 41748
rect 11900 41970 11956 41972
rect 11900 41918 11902 41970
rect 11902 41918 11954 41970
rect 11954 41918 11956 41970
rect 11900 41916 11956 41918
rect 11676 41468 11732 41524
rect 12460 41468 12516 41524
rect 11900 41410 11956 41412
rect 11900 41358 11902 41410
rect 11902 41358 11954 41410
rect 11954 41358 11956 41410
rect 11900 41356 11956 41358
rect 12012 41186 12068 41188
rect 12012 41134 12014 41186
rect 12014 41134 12066 41186
rect 12066 41134 12068 41186
rect 12012 41132 12068 41134
rect 12572 41186 12628 41188
rect 12572 41134 12574 41186
rect 12574 41134 12626 41186
rect 12626 41134 12628 41186
rect 12572 41132 12628 41134
rect 11900 41074 11956 41076
rect 11900 41022 11902 41074
rect 11902 41022 11954 41074
rect 11954 41022 11956 41074
rect 11900 41020 11956 41022
rect 12460 40572 12516 40628
rect 13580 42642 13636 42644
rect 13580 42590 13582 42642
rect 13582 42590 13634 42642
rect 13634 42590 13636 42642
rect 13580 42588 13636 42590
rect 13580 41804 13636 41860
rect 13020 41132 13076 41188
rect 13692 40572 13748 40628
rect 13804 40796 13860 40852
rect 13356 40402 13412 40404
rect 13356 40350 13358 40402
rect 13358 40350 13410 40402
rect 13410 40350 13412 40402
rect 13356 40348 13412 40350
rect 13916 40402 13972 40404
rect 13916 40350 13918 40402
rect 13918 40350 13970 40402
rect 13970 40350 13972 40402
rect 13916 40348 13972 40350
rect 11676 38780 11732 38836
rect 11452 36876 11508 36932
rect 10220 31276 10276 31332
rect 10892 36204 10948 36260
rect 10444 33122 10500 33124
rect 10444 33070 10446 33122
rect 10446 33070 10498 33122
rect 10498 33070 10500 33122
rect 10444 33068 10500 33070
rect 10444 32060 10500 32116
rect 10556 32284 10612 32340
rect 9436 31218 9492 31220
rect 9436 31166 9438 31218
rect 9438 31166 9490 31218
rect 9490 31166 9492 31218
rect 9436 31164 9492 31166
rect 9884 31164 9940 31220
rect 9212 30268 9268 30324
rect 9772 30994 9828 30996
rect 9772 30942 9774 30994
rect 9774 30942 9826 30994
rect 9826 30942 9828 30994
rect 9772 30940 9828 30942
rect 9772 30268 9828 30324
rect 8876 29932 8932 29988
rect 8988 28812 9044 28868
rect 9100 28642 9156 28644
rect 9100 28590 9102 28642
rect 9102 28590 9154 28642
rect 9154 28590 9156 28642
rect 9100 28588 9156 28590
rect 8988 28476 9044 28532
rect 8092 27970 8148 27972
rect 8092 27918 8094 27970
rect 8094 27918 8146 27970
rect 8146 27918 8148 27970
rect 8092 27916 8148 27918
rect 9548 28812 9604 28868
rect 9324 28642 9380 28644
rect 9324 28590 9326 28642
rect 9326 28590 9378 28642
rect 9378 28590 9380 28642
rect 9324 28588 9380 28590
rect 9996 30994 10052 30996
rect 9996 30942 9998 30994
rect 9998 30942 10050 30994
rect 10050 30942 10052 30994
rect 9996 30940 10052 30942
rect 10668 31948 10724 32004
rect 11228 36092 11284 36148
rect 11004 32562 11060 32564
rect 11004 32510 11006 32562
rect 11006 32510 11058 32562
rect 11058 32510 11060 32562
rect 11004 32508 11060 32510
rect 10780 31890 10836 31892
rect 10780 31838 10782 31890
rect 10782 31838 10834 31890
rect 10834 31838 10836 31890
rect 10780 31836 10836 31838
rect 11228 31388 11284 31444
rect 10892 30940 10948 30996
rect 10220 30268 10276 30324
rect 10332 30156 10388 30212
rect 10220 29484 10276 29540
rect 9996 28588 10052 28644
rect 9436 28082 9492 28084
rect 9436 28030 9438 28082
rect 9438 28030 9490 28082
rect 9490 28030 9492 28082
rect 9436 28028 9492 28030
rect 9548 27970 9604 27972
rect 9548 27918 9550 27970
rect 9550 27918 9602 27970
rect 9602 27918 9604 27970
rect 9548 27916 9604 27918
rect 8204 27580 8260 27636
rect 8316 27244 8372 27300
rect 8540 27634 8596 27636
rect 8540 27582 8542 27634
rect 8542 27582 8594 27634
rect 8594 27582 8596 27634
rect 8540 27580 8596 27582
rect 7420 25788 7476 25844
rect 6860 25730 6916 25732
rect 6860 25678 6862 25730
rect 6862 25678 6914 25730
rect 6914 25678 6916 25730
rect 6860 25676 6916 25678
rect 6748 23884 6804 23940
rect 8764 26684 8820 26740
rect 8876 27804 8932 27860
rect 9436 27804 9492 27860
rect 9100 26796 9156 26852
rect 8092 26178 8148 26180
rect 8092 26126 8094 26178
rect 8094 26126 8146 26178
rect 8146 26126 8148 26178
rect 8092 26124 8148 26126
rect 7980 25788 8036 25844
rect 8204 25676 8260 25732
rect 8428 26012 8484 26068
rect 7756 25116 7812 25172
rect 7644 24050 7700 24052
rect 7644 23998 7646 24050
rect 7646 23998 7698 24050
rect 7698 23998 7700 24050
rect 7644 23996 7700 23998
rect 6300 22988 6356 23044
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4284 20802 4340 20804
rect 4284 20750 4286 20802
rect 4286 20750 4338 20802
rect 4338 20750 4340 20802
rect 4284 20748 4340 20750
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5068 17778 5124 17780
rect 5068 17726 5070 17778
rect 5070 17726 5122 17778
rect 5122 17726 5124 17778
rect 5068 17724 5124 17726
rect 3948 17164 4004 17220
rect 5852 20748 5908 20804
rect 6636 22204 6692 22260
rect 6524 18450 6580 18452
rect 6524 18398 6526 18450
rect 6526 18398 6578 18450
rect 6578 18398 6580 18450
rect 6524 18396 6580 18398
rect 4060 16994 4116 16996
rect 4060 16942 4062 16994
rect 4062 16942 4114 16994
rect 4114 16942 4116 16994
rect 4060 16940 4116 16942
rect 3500 16492 3556 16548
rect 5740 16828 5796 16884
rect 3164 15426 3220 15428
rect 3164 15374 3166 15426
rect 3166 15374 3218 15426
rect 3218 15374 3220 15426
rect 3164 15372 3220 15374
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 5740 16210 5796 16212
rect 5740 16158 5742 16210
rect 5742 16158 5794 16210
rect 5794 16158 5796 16210
rect 5740 16156 5796 16158
rect 5292 15202 5348 15204
rect 5292 15150 5294 15202
rect 5294 15150 5346 15202
rect 5346 15150 5348 15202
rect 5292 15148 5348 15150
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3500 13692 3556 13748
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 7420 23548 7476 23604
rect 7308 23154 7364 23156
rect 7308 23102 7310 23154
rect 7310 23102 7362 23154
rect 7362 23102 7364 23154
rect 7308 23100 7364 23102
rect 6188 17724 6244 17780
rect 7084 22764 7140 22820
rect 6076 16828 6132 16884
rect 6188 16770 6244 16772
rect 6188 16718 6190 16770
rect 6190 16718 6242 16770
rect 6242 16718 6244 16770
rect 6188 16716 6244 16718
rect 5964 15932 6020 15988
rect 6748 17554 6804 17556
rect 6748 17502 6750 17554
rect 6750 17502 6802 17554
rect 6802 17502 6804 17554
rect 6748 17500 6804 17502
rect 6972 17554 7028 17556
rect 6972 17502 6974 17554
rect 6974 17502 7026 17554
rect 7026 17502 7028 17554
rect 6972 17500 7028 17502
rect 7196 22428 7252 22484
rect 8204 24780 8260 24836
rect 7868 23938 7924 23940
rect 7868 23886 7870 23938
rect 7870 23886 7922 23938
rect 7922 23886 7924 23938
rect 7868 23884 7924 23886
rect 7756 22988 7812 23044
rect 7644 22540 7700 22596
rect 7532 22092 7588 22148
rect 7644 21474 7700 21476
rect 7644 21422 7646 21474
rect 7646 21422 7698 21474
rect 7698 21422 7700 21474
rect 7644 21420 7700 21422
rect 7196 19068 7252 19124
rect 7196 18450 7252 18452
rect 7196 18398 7198 18450
rect 7198 18398 7250 18450
rect 7250 18398 7252 18450
rect 7196 18396 7252 18398
rect 7980 23154 8036 23156
rect 7980 23102 7982 23154
rect 7982 23102 8034 23154
rect 8034 23102 8036 23154
rect 7980 23100 8036 23102
rect 8316 23042 8372 23044
rect 8316 22990 8318 23042
rect 8318 22990 8370 23042
rect 8370 22990 8372 23042
rect 8316 22988 8372 22990
rect 8316 22146 8372 22148
rect 8316 22094 8318 22146
rect 8318 22094 8370 22146
rect 8370 22094 8372 22146
rect 8316 22092 8372 22094
rect 8652 25228 8708 25284
rect 8988 24780 9044 24836
rect 8876 24444 8932 24500
rect 8764 23996 8820 24052
rect 8764 22258 8820 22260
rect 8764 22206 8766 22258
rect 8766 22206 8818 22258
rect 8818 22206 8820 22258
rect 8764 22204 8820 22206
rect 9772 27746 9828 27748
rect 9772 27694 9774 27746
rect 9774 27694 9826 27746
rect 9826 27694 9828 27746
rect 9772 27692 9828 27694
rect 9884 27580 9940 27636
rect 11564 36764 11620 36820
rect 11900 38722 11956 38724
rect 11900 38670 11902 38722
rect 11902 38670 11954 38722
rect 11954 38670 11956 38722
rect 11900 38668 11956 38670
rect 11900 38444 11956 38500
rect 12572 39058 12628 39060
rect 12572 39006 12574 39058
rect 12574 39006 12626 39058
rect 12626 39006 12628 39058
rect 12572 39004 12628 39006
rect 12460 38892 12516 38948
rect 12124 38834 12180 38836
rect 12124 38782 12126 38834
rect 12126 38782 12178 38834
rect 12178 38782 12180 38834
rect 12124 38780 12180 38782
rect 12460 38444 12516 38500
rect 12460 37378 12516 37380
rect 12460 37326 12462 37378
rect 12462 37326 12514 37378
rect 12514 37326 12516 37378
rect 12460 37324 12516 37326
rect 12796 37324 12852 37380
rect 12012 37212 12068 37268
rect 12572 37212 12628 37268
rect 12012 36706 12068 36708
rect 12012 36654 12014 36706
rect 12014 36654 12066 36706
rect 12066 36654 12068 36706
rect 12012 36652 12068 36654
rect 12236 36594 12292 36596
rect 12236 36542 12238 36594
rect 12238 36542 12290 36594
rect 12290 36542 12292 36594
rect 12236 36540 12292 36542
rect 12460 36988 12516 37044
rect 11788 36370 11844 36372
rect 11788 36318 11790 36370
rect 11790 36318 11842 36370
rect 11842 36318 11844 36370
rect 11788 36316 11844 36318
rect 11676 36092 11732 36148
rect 11564 35980 11620 36036
rect 11676 35868 11732 35924
rect 12124 35084 12180 35140
rect 11788 34524 11844 34580
rect 12236 36092 12292 36148
rect 12460 36092 12516 36148
rect 12684 37100 12740 37156
rect 12908 36428 12964 36484
rect 12684 36316 12740 36372
rect 12348 35308 12404 35364
rect 12236 34524 12292 34580
rect 12572 34802 12628 34804
rect 12572 34750 12574 34802
rect 12574 34750 12626 34802
rect 12626 34750 12628 34802
rect 12572 34748 12628 34750
rect 12908 34748 12964 34804
rect 12012 33404 12068 33460
rect 11564 31164 11620 31220
rect 12348 32620 12404 32676
rect 12684 34300 12740 34356
rect 12796 33292 12852 33348
rect 12684 32620 12740 32676
rect 11452 31052 11508 31108
rect 12124 31778 12180 31780
rect 12124 31726 12126 31778
rect 12126 31726 12178 31778
rect 12178 31726 12180 31778
rect 12124 31724 12180 31726
rect 11900 30940 11956 30996
rect 11788 30156 11844 30212
rect 11340 30044 11396 30100
rect 11788 29484 11844 29540
rect 11340 28476 11396 28532
rect 9996 27020 10052 27076
rect 11564 27356 11620 27412
rect 10444 27074 10500 27076
rect 10444 27022 10446 27074
rect 10446 27022 10498 27074
rect 10498 27022 10500 27074
rect 10444 27020 10500 27022
rect 10220 26796 10276 26852
rect 9996 26012 10052 26068
rect 9772 23996 9828 24052
rect 9884 24556 9940 24612
rect 9436 22764 9492 22820
rect 9100 22652 9156 22708
rect 10668 26012 10724 26068
rect 10668 23884 10724 23940
rect 9996 22204 10052 22260
rect 8428 21420 8484 21476
rect 8316 20524 8372 20580
rect 7980 19906 8036 19908
rect 7980 19854 7982 19906
rect 7982 19854 8034 19906
rect 8034 19854 8036 19906
rect 7980 19852 8036 19854
rect 8428 19628 8484 19684
rect 8316 19180 8372 19236
rect 8988 21698 9044 21700
rect 8988 21646 8990 21698
rect 8990 21646 9042 21698
rect 9042 21646 9044 21698
rect 8988 21644 9044 21646
rect 8988 21196 9044 21252
rect 9100 20578 9156 20580
rect 9100 20526 9102 20578
rect 9102 20526 9154 20578
rect 9154 20526 9156 20578
rect 9100 20524 9156 20526
rect 9660 21586 9716 21588
rect 9660 21534 9662 21586
rect 9662 21534 9714 21586
rect 9714 21534 9716 21586
rect 9660 21532 9716 21534
rect 10108 21980 10164 22036
rect 10108 21532 10164 21588
rect 10668 21532 10724 21588
rect 12460 32508 12516 32564
rect 12908 32562 12964 32564
rect 12908 32510 12910 32562
rect 12910 32510 12962 32562
rect 12962 32510 12964 32562
rect 12908 32508 12964 32510
rect 12684 31500 12740 31556
rect 13916 39900 13972 39956
rect 13692 39564 13748 39620
rect 13468 38892 13524 38948
rect 13916 39058 13972 39060
rect 13916 39006 13918 39058
rect 13918 39006 13970 39058
rect 13970 39006 13972 39058
rect 13916 39004 13972 39006
rect 13692 38780 13748 38836
rect 13244 37154 13300 37156
rect 13244 37102 13246 37154
rect 13246 37102 13298 37154
rect 13298 37102 13300 37154
rect 13244 37100 13300 37102
rect 13356 36652 13412 36708
rect 13132 36540 13188 36596
rect 13132 35308 13188 35364
rect 13916 37996 13972 38052
rect 13804 37490 13860 37492
rect 13804 37438 13806 37490
rect 13806 37438 13858 37490
rect 13858 37438 13860 37490
rect 13804 37436 13860 37438
rect 15260 45612 15316 45668
rect 14700 45164 14756 45220
rect 14812 44098 14868 44100
rect 14812 44046 14814 44098
rect 14814 44046 14866 44098
rect 14866 44046 14868 44098
rect 14812 44044 14868 44046
rect 15148 44098 15204 44100
rect 15148 44046 15150 44098
rect 15150 44046 15202 44098
rect 15202 44046 15204 44098
rect 15148 44044 15204 44046
rect 14252 43596 14308 43652
rect 14812 43426 14868 43428
rect 14812 43374 14814 43426
rect 14814 43374 14866 43426
rect 14866 43374 14868 43426
rect 14812 43372 14868 43374
rect 14700 42028 14756 42084
rect 14364 40796 14420 40852
rect 14140 39394 14196 39396
rect 14140 39342 14142 39394
rect 14142 39342 14194 39394
rect 14194 39342 14196 39394
rect 14140 39340 14196 39342
rect 14252 39228 14308 39284
rect 14364 39116 14420 39172
rect 15036 42028 15092 42084
rect 15036 39730 15092 39732
rect 15036 39678 15038 39730
rect 15038 39678 15090 39730
rect 15090 39678 15092 39730
rect 15036 39676 15092 39678
rect 16380 43596 16436 43652
rect 15484 42476 15540 42532
rect 14700 39116 14756 39172
rect 14588 38780 14644 38836
rect 14700 38668 14756 38724
rect 14364 38332 14420 38388
rect 15036 38780 15092 38836
rect 18956 45724 19012 45780
rect 17948 43650 18004 43652
rect 17948 43598 17950 43650
rect 17950 43598 18002 43650
rect 18002 43598 18004 43650
rect 17948 43596 18004 43598
rect 17276 42812 17332 42868
rect 16380 42476 16436 42532
rect 16604 42588 16660 42644
rect 16380 40348 16436 40404
rect 15708 39730 15764 39732
rect 15708 39678 15710 39730
rect 15710 39678 15762 39730
rect 15762 39678 15764 39730
rect 15708 39676 15764 39678
rect 14028 36876 14084 36932
rect 13580 36594 13636 36596
rect 13580 36542 13582 36594
rect 13582 36542 13634 36594
rect 13634 36542 13636 36594
rect 13580 36540 13636 36542
rect 13468 36482 13524 36484
rect 13468 36430 13470 36482
rect 13470 36430 13522 36482
rect 13522 36430 13524 36482
rect 13468 36428 13524 36430
rect 14028 36540 14084 36596
rect 13468 36204 13524 36260
rect 13916 36204 13972 36260
rect 13356 35532 13412 35588
rect 13132 34354 13188 34356
rect 13132 34302 13134 34354
rect 13134 34302 13186 34354
rect 13186 34302 13188 34354
rect 13132 34300 13188 34302
rect 14028 35084 14084 35140
rect 13692 35026 13748 35028
rect 13692 34974 13694 35026
rect 13694 34974 13746 35026
rect 13746 34974 13748 35026
rect 13692 34972 13748 34974
rect 13468 34860 13524 34916
rect 13356 31724 13412 31780
rect 13692 32620 13748 32676
rect 13468 31500 13524 31556
rect 13468 30492 13524 30548
rect 13244 30380 13300 30436
rect 13580 30380 13636 30436
rect 14364 35698 14420 35700
rect 14364 35646 14366 35698
rect 14366 35646 14418 35698
rect 14418 35646 14420 35698
rect 14364 35644 14420 35646
rect 15148 37100 15204 37156
rect 14812 36876 14868 36932
rect 14812 36428 14868 36484
rect 14700 35868 14756 35924
rect 14812 36204 14868 36260
rect 14476 34524 14532 34580
rect 14364 32562 14420 32564
rect 14364 32510 14366 32562
rect 14366 32510 14418 32562
rect 14418 32510 14420 32562
rect 14364 32508 14420 32510
rect 15596 36594 15652 36596
rect 15596 36542 15598 36594
rect 15598 36542 15650 36594
rect 15650 36542 15652 36594
rect 15596 36540 15652 36542
rect 13916 31836 13972 31892
rect 14028 31724 14084 31780
rect 13020 30156 13076 30212
rect 13804 31612 13860 31668
rect 12348 29484 12404 29540
rect 13132 30044 13188 30100
rect 13692 29538 13748 29540
rect 13692 29486 13694 29538
rect 13694 29486 13746 29538
rect 13746 29486 13748 29538
rect 13692 29484 13748 29486
rect 15036 35868 15092 35924
rect 14588 31218 14644 31220
rect 14588 31166 14590 31218
rect 14590 31166 14642 31218
rect 14642 31166 14644 31218
rect 14588 31164 14644 31166
rect 14252 30882 14308 30884
rect 14252 30830 14254 30882
rect 14254 30830 14306 30882
rect 14306 30830 14308 30882
rect 14252 30828 14308 30830
rect 14476 30828 14532 30884
rect 14812 30770 14868 30772
rect 14812 30718 14814 30770
rect 14814 30718 14866 30770
rect 14866 30718 14868 30770
rect 14812 30716 14868 30718
rect 14028 30492 14084 30548
rect 13916 30268 13972 30324
rect 15036 30380 15092 30436
rect 15484 36428 15540 36484
rect 15484 36204 15540 36260
rect 16044 39676 16100 39732
rect 16156 39340 16212 39396
rect 16268 39116 16324 39172
rect 16492 39004 16548 39060
rect 15820 37266 15876 37268
rect 15820 37214 15822 37266
rect 15822 37214 15874 37266
rect 15874 37214 15876 37266
rect 15820 37212 15876 37214
rect 16156 36540 16212 36596
rect 15708 35922 15764 35924
rect 15708 35870 15710 35922
rect 15710 35870 15762 35922
rect 15762 35870 15764 35922
rect 15708 35868 15764 35870
rect 16044 36204 16100 36260
rect 15932 35196 15988 35252
rect 15372 34524 15428 34580
rect 15260 31106 15316 31108
rect 15260 31054 15262 31106
rect 15262 31054 15314 31106
rect 15314 31054 15316 31106
rect 15260 31052 15316 31054
rect 15596 32508 15652 32564
rect 14252 30210 14308 30212
rect 14252 30158 14254 30210
rect 14254 30158 14306 30210
rect 14306 30158 14308 30210
rect 14252 30156 14308 30158
rect 14700 30210 14756 30212
rect 14700 30158 14702 30210
rect 14702 30158 14754 30210
rect 14754 30158 14756 30210
rect 14700 30156 14756 30158
rect 15036 30156 15092 30212
rect 14476 29986 14532 29988
rect 14476 29934 14478 29986
rect 14478 29934 14530 29986
rect 14530 29934 14532 29986
rect 14476 29932 14532 29934
rect 14812 29820 14868 29876
rect 13132 28364 13188 28420
rect 13692 28252 13748 28308
rect 12012 25564 12068 25620
rect 13020 26460 13076 26516
rect 11116 24668 11172 24724
rect 11788 24722 11844 24724
rect 11788 24670 11790 24722
rect 11790 24670 11842 24722
rect 11842 24670 11844 24722
rect 11788 24668 11844 24670
rect 12236 24668 12292 24724
rect 11676 24444 11732 24500
rect 11676 23772 11732 23828
rect 11452 21810 11508 21812
rect 11452 21758 11454 21810
rect 11454 21758 11506 21810
rect 11506 21758 11508 21810
rect 11452 21756 11508 21758
rect 12796 24722 12852 24724
rect 12796 24670 12798 24722
rect 12798 24670 12850 24722
rect 12850 24670 12852 24722
rect 12796 24668 12852 24670
rect 12460 24108 12516 24164
rect 11900 23772 11956 23828
rect 12684 23826 12740 23828
rect 12684 23774 12686 23826
rect 12686 23774 12738 23826
rect 12738 23774 12740 23826
rect 12684 23772 12740 23774
rect 12684 23548 12740 23604
rect 12236 23042 12292 23044
rect 12236 22990 12238 23042
rect 12238 22990 12290 23042
rect 12290 22990 12292 23042
rect 12236 22988 12292 22990
rect 11564 21644 11620 21700
rect 11900 21868 11956 21924
rect 10892 20914 10948 20916
rect 10892 20862 10894 20914
rect 10894 20862 10946 20914
rect 10946 20862 10948 20914
rect 10892 20860 10948 20862
rect 9436 20578 9492 20580
rect 9436 20526 9438 20578
rect 9438 20526 9490 20578
rect 9490 20526 9492 20578
rect 9436 20524 9492 20526
rect 9996 20412 10052 20468
rect 8764 19852 8820 19908
rect 9660 19628 9716 19684
rect 8876 19010 8932 19012
rect 8876 18958 8878 19010
rect 8878 18958 8930 19010
rect 8930 18958 8932 19010
rect 8876 18956 8932 18958
rect 9772 19234 9828 19236
rect 9772 19182 9774 19234
rect 9774 19182 9826 19234
rect 9826 19182 9828 19234
rect 9772 19180 9828 19182
rect 9660 18620 9716 18676
rect 8876 18508 8932 18564
rect 8652 17836 8708 17892
rect 6748 17052 6804 17108
rect 6860 16994 6916 16996
rect 6860 16942 6862 16994
rect 6862 16942 6914 16994
rect 6914 16942 6916 16994
rect 6860 16940 6916 16942
rect 7084 16994 7140 16996
rect 7084 16942 7086 16994
rect 7086 16942 7138 16994
rect 7138 16942 7140 16994
rect 7084 16940 7140 16942
rect 7420 17052 7476 17108
rect 8204 17388 8260 17444
rect 6188 15484 6244 15540
rect 6972 16098 7028 16100
rect 6972 16046 6974 16098
rect 6974 16046 7026 16098
rect 7026 16046 7028 16098
rect 6972 16044 7028 16046
rect 6860 15538 6916 15540
rect 6860 15486 6862 15538
rect 6862 15486 6914 15538
rect 6914 15486 6916 15538
rect 6860 15484 6916 15486
rect 7084 15932 7140 15988
rect 6748 15372 6804 15428
rect 6300 15148 6356 15204
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5516 14476 5572 14532
rect 3052 10668 3108 10724
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 2492 4226 2548 4228
rect 2492 4174 2494 4226
rect 2494 4174 2546 4226
rect 2546 4174 2548 4226
rect 2492 4172 2548 4174
rect 1708 3276 1764 3332
rect 1708 2044 1764 2100
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 6076 11676 6132 11732
rect 5516 9212 5572 9268
rect 7196 15820 7252 15876
rect 7420 16716 7476 16772
rect 7868 16882 7924 16884
rect 7868 16830 7870 16882
rect 7870 16830 7922 16882
rect 7922 16830 7924 16882
rect 7868 16828 7924 16830
rect 7756 16716 7812 16772
rect 8204 16716 8260 16772
rect 7868 16098 7924 16100
rect 7868 16046 7870 16098
rect 7870 16046 7922 16098
rect 7922 16046 7924 16098
rect 7868 16044 7924 16046
rect 8092 15986 8148 15988
rect 8092 15934 8094 15986
rect 8094 15934 8146 15986
rect 8146 15934 8148 15986
rect 8092 15932 8148 15934
rect 7644 15874 7700 15876
rect 7644 15822 7646 15874
rect 7646 15822 7698 15874
rect 7698 15822 7700 15874
rect 7644 15820 7700 15822
rect 7756 15538 7812 15540
rect 7756 15486 7758 15538
rect 7758 15486 7810 15538
rect 7810 15486 7812 15538
rect 7756 15484 7812 15486
rect 8204 13580 8260 13636
rect 2940 3276 2996 3332
rect 8428 17554 8484 17556
rect 8428 17502 8430 17554
rect 8430 17502 8482 17554
rect 8482 17502 8484 17554
rect 8428 17500 8484 17502
rect 8540 17388 8596 17444
rect 8764 16716 8820 16772
rect 8652 15986 8708 15988
rect 8652 15934 8654 15986
rect 8654 15934 8706 15986
rect 8706 15934 8708 15986
rect 8652 15932 8708 15934
rect 9772 18562 9828 18564
rect 9772 18510 9774 18562
rect 9774 18510 9826 18562
rect 9826 18510 9828 18562
rect 9772 18508 9828 18510
rect 9772 17948 9828 18004
rect 9100 17836 9156 17892
rect 8988 16940 9044 16996
rect 9324 16716 9380 16772
rect 9772 16828 9828 16884
rect 11004 19964 11060 20020
rect 10668 19906 10724 19908
rect 10668 19854 10670 19906
rect 10670 19854 10722 19906
rect 10722 19854 10724 19906
rect 10668 19852 10724 19854
rect 10668 19346 10724 19348
rect 10668 19294 10670 19346
rect 10670 19294 10722 19346
rect 10722 19294 10724 19346
rect 10668 19292 10724 19294
rect 10108 18508 10164 18564
rect 11004 18956 11060 19012
rect 10668 18508 10724 18564
rect 11004 17276 11060 17332
rect 10556 16268 10612 16324
rect 10668 16716 10724 16772
rect 9548 15538 9604 15540
rect 9548 15486 9550 15538
rect 9550 15486 9602 15538
rect 9602 15486 9604 15538
rect 9548 15484 9604 15486
rect 8428 14140 8484 14196
rect 9660 13634 9716 13636
rect 9660 13582 9662 13634
rect 9662 13582 9714 13634
rect 9714 13582 9716 13634
rect 9660 13580 9716 13582
rect 9996 15484 10052 15540
rect 9884 14140 9940 14196
rect 10332 15148 10388 15204
rect 10892 15202 10948 15204
rect 10892 15150 10894 15202
rect 10894 15150 10946 15202
rect 10946 15150 10948 15202
rect 10892 15148 10948 15150
rect 11564 19964 11620 20020
rect 11340 19516 11396 19572
rect 12012 22092 12068 22148
rect 12236 21756 12292 21812
rect 12124 21586 12180 21588
rect 12124 21534 12126 21586
rect 12126 21534 12178 21586
rect 12178 21534 12180 21586
rect 12124 21532 12180 21534
rect 11900 19906 11956 19908
rect 11900 19854 11902 19906
rect 11902 19854 11954 19906
rect 11954 19854 11956 19906
rect 11900 19852 11956 19854
rect 11900 19516 11956 19572
rect 11564 18562 11620 18564
rect 11564 18510 11566 18562
rect 11566 18510 11618 18562
rect 11618 18510 11620 18562
rect 11564 18508 11620 18510
rect 12572 21196 12628 21252
rect 12348 20914 12404 20916
rect 12348 20862 12350 20914
rect 12350 20862 12402 20914
rect 12402 20862 12404 20914
rect 12348 20860 12404 20862
rect 13580 24108 13636 24164
rect 13580 23772 13636 23828
rect 13580 23212 13636 23268
rect 13580 22258 13636 22260
rect 13580 22206 13582 22258
rect 13582 22206 13634 22258
rect 13634 22206 13636 22258
rect 13580 22204 13636 22206
rect 13468 21756 13524 21812
rect 14028 28364 14084 28420
rect 14028 26236 14084 26292
rect 13916 25340 13972 25396
rect 13916 24780 13972 24836
rect 14028 23826 14084 23828
rect 14028 23774 14030 23826
rect 14030 23774 14082 23826
rect 14082 23774 14084 23826
rect 14028 23772 14084 23774
rect 14028 22988 14084 23044
rect 14028 22370 14084 22372
rect 14028 22318 14030 22370
rect 14030 22318 14082 22370
rect 14082 22318 14084 22370
rect 14028 22316 14084 22318
rect 13804 22146 13860 22148
rect 13804 22094 13806 22146
rect 13806 22094 13858 22146
rect 13858 22094 13860 22146
rect 13804 22092 13860 22094
rect 12908 21026 12964 21028
rect 12908 20974 12910 21026
rect 12910 20974 12962 21026
rect 12962 20974 12964 21026
rect 12908 20972 12964 20974
rect 12796 20860 12852 20916
rect 12348 19628 12404 19684
rect 13804 20076 13860 20132
rect 12908 19852 12964 19908
rect 12796 19516 12852 19572
rect 12572 19404 12628 19460
rect 12348 19346 12404 19348
rect 12348 19294 12350 19346
rect 12350 19294 12402 19346
rect 12402 19294 12404 19346
rect 12348 19292 12404 19294
rect 13804 19628 13860 19684
rect 14364 26850 14420 26852
rect 14364 26798 14366 26850
rect 14366 26798 14418 26850
rect 14418 26798 14420 26850
rect 14364 26796 14420 26798
rect 14252 25394 14308 25396
rect 14252 25342 14254 25394
rect 14254 25342 14306 25394
rect 14306 25342 14308 25394
rect 14252 25340 14308 25342
rect 15148 30044 15204 30100
rect 14812 27858 14868 27860
rect 14812 27806 14814 27858
rect 14814 27806 14866 27858
rect 14866 27806 14868 27858
rect 14812 27804 14868 27806
rect 15036 28364 15092 28420
rect 16044 31276 16100 31332
rect 15708 30098 15764 30100
rect 15708 30046 15710 30098
rect 15710 30046 15762 30098
rect 15762 30046 15764 30098
rect 15708 30044 15764 30046
rect 16044 30380 16100 30436
rect 16156 30492 16212 30548
rect 15932 30156 15988 30212
rect 16940 42140 16996 42196
rect 16828 40460 16884 40516
rect 16828 39730 16884 39732
rect 16828 39678 16830 39730
rect 16830 39678 16882 39730
rect 16882 39678 16884 39730
rect 16828 39676 16884 39678
rect 16716 39340 16772 39396
rect 16604 36876 16660 36932
rect 16380 36092 16436 36148
rect 16716 34076 16772 34132
rect 16828 35308 16884 35364
rect 17388 42140 17444 42196
rect 17836 42588 17892 42644
rect 18172 43260 18228 43316
rect 18284 45388 18340 45444
rect 18060 42924 18116 42980
rect 18172 41074 18228 41076
rect 18172 41022 18174 41074
rect 18174 41022 18226 41074
rect 18226 41022 18228 41074
rect 18172 41020 18228 41022
rect 17724 40684 17780 40740
rect 17388 39004 17444 39060
rect 17052 38556 17108 38612
rect 17836 38780 17892 38836
rect 17164 36540 17220 36596
rect 17612 38332 17668 38388
rect 18060 40348 18116 40404
rect 18060 39116 18116 39172
rect 18508 43596 18564 43652
rect 18732 43260 18788 43316
rect 18508 42588 18564 42644
rect 18396 42476 18452 42532
rect 18508 42140 18564 42196
rect 18396 42082 18452 42084
rect 18396 42030 18398 42082
rect 18398 42030 18450 42082
rect 18450 42030 18452 42082
rect 18396 42028 18452 42030
rect 18060 37378 18116 37380
rect 18060 37326 18062 37378
rect 18062 37326 18114 37378
rect 18114 37326 18116 37378
rect 18060 37324 18116 37326
rect 18396 41804 18452 41860
rect 17500 35420 17556 35476
rect 17388 35308 17444 35364
rect 17948 36204 18004 36260
rect 18060 35756 18116 35812
rect 18844 42252 18900 42308
rect 18732 41804 18788 41860
rect 18844 42028 18900 42084
rect 18508 41132 18564 41188
rect 18732 41074 18788 41076
rect 18732 41022 18734 41074
rect 18734 41022 18786 41074
rect 18786 41022 18788 41074
rect 18732 41020 18788 41022
rect 18620 40684 18676 40740
rect 18508 40572 18564 40628
rect 18620 38780 18676 38836
rect 18508 38668 18564 38724
rect 18844 38946 18900 38948
rect 18844 38894 18846 38946
rect 18846 38894 18898 38946
rect 18898 38894 18900 38946
rect 18844 38892 18900 38894
rect 18732 37772 18788 37828
rect 18508 36988 18564 37044
rect 18284 35420 18340 35476
rect 18060 35308 18116 35364
rect 18620 36092 18676 36148
rect 18620 35420 18676 35476
rect 18844 37100 18900 37156
rect 19068 45388 19124 45444
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19180 43596 19236 43652
rect 20412 43426 20468 43428
rect 20412 43374 20414 43426
rect 20414 43374 20466 43426
rect 20466 43374 20468 43426
rect 20412 43372 20468 43374
rect 19404 43314 19460 43316
rect 19404 43262 19406 43314
rect 19406 43262 19458 43314
rect 19458 43262 19460 43314
rect 19404 43260 19460 43262
rect 20636 43148 20692 43204
rect 19740 42812 19796 42868
rect 19404 42252 19460 42308
rect 19516 42476 19572 42532
rect 19516 42028 19572 42084
rect 19404 41916 19460 41972
rect 19292 40348 19348 40404
rect 19180 38722 19236 38724
rect 19180 38670 19182 38722
rect 19182 38670 19234 38722
rect 19234 38670 19236 38722
rect 19180 38668 19236 38670
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19404 38108 19460 38164
rect 20076 42140 20132 42196
rect 24108 45836 24164 45892
rect 21756 45724 21812 45780
rect 23100 45666 23156 45668
rect 23100 45614 23102 45666
rect 23102 45614 23154 45666
rect 23154 45614 23156 45666
rect 23100 45612 23156 45614
rect 22764 44268 22820 44324
rect 20972 44156 21028 44212
rect 22428 44210 22484 44212
rect 22428 44158 22430 44210
rect 22430 44158 22482 44210
rect 22482 44158 22484 44210
rect 22428 44156 22484 44158
rect 21308 43596 21364 43652
rect 21868 43596 21924 43652
rect 21532 43372 21588 43428
rect 21420 43036 21476 43092
rect 20748 41916 20804 41972
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20412 41020 20468 41076
rect 20300 39452 20356 39508
rect 19628 39340 19684 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20636 39340 20692 39396
rect 21308 39394 21364 39396
rect 21308 39342 21310 39394
rect 21310 39342 21362 39394
rect 21362 39342 21364 39394
rect 21308 39340 21364 39342
rect 20300 38892 20356 38948
rect 20300 37826 20356 37828
rect 20300 37774 20302 37826
rect 20302 37774 20354 37826
rect 20354 37774 20356 37826
rect 20300 37772 20356 37774
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20524 37324 20580 37380
rect 19068 37154 19124 37156
rect 19068 37102 19070 37154
rect 19070 37102 19122 37154
rect 19122 37102 19124 37154
rect 19068 37100 19124 37102
rect 19292 37042 19348 37044
rect 19292 36990 19294 37042
rect 19294 36990 19346 37042
rect 19346 36990 19348 37042
rect 19292 36988 19348 36990
rect 19292 36428 19348 36484
rect 18844 36258 18900 36260
rect 18844 36206 18846 36258
rect 18846 36206 18898 36258
rect 18898 36206 18900 36258
rect 18844 36204 18900 36206
rect 19180 36316 19236 36372
rect 18844 35756 18900 35812
rect 19292 35810 19348 35812
rect 19292 35758 19294 35810
rect 19294 35758 19346 35810
rect 19346 35758 19348 35810
rect 19292 35756 19348 35758
rect 18844 35586 18900 35588
rect 18844 35534 18846 35586
rect 18846 35534 18898 35586
rect 18898 35534 18900 35586
rect 18844 35532 18900 35534
rect 18732 34636 18788 34692
rect 17724 33458 17780 33460
rect 17724 33406 17726 33458
rect 17726 33406 17778 33458
rect 17778 33406 17780 33458
rect 17724 33404 17780 33406
rect 17836 33346 17892 33348
rect 17836 33294 17838 33346
rect 17838 33294 17890 33346
rect 17890 33294 17892 33346
rect 17836 33292 17892 33294
rect 17052 33234 17108 33236
rect 17052 33182 17054 33234
rect 17054 33182 17106 33234
rect 17106 33182 17108 33234
rect 17052 33180 17108 33182
rect 16716 30210 16772 30212
rect 16716 30158 16718 30210
rect 16718 30158 16770 30210
rect 16770 30158 16772 30210
rect 16716 30156 16772 30158
rect 16044 29650 16100 29652
rect 16044 29598 16046 29650
rect 16046 29598 16098 29650
rect 16098 29598 16100 29650
rect 16044 29596 16100 29598
rect 16380 29708 16436 29764
rect 15820 29372 15876 29428
rect 15484 28642 15540 28644
rect 15484 28590 15486 28642
rect 15486 28590 15538 28642
rect 15538 28590 15540 28642
rect 15484 28588 15540 28590
rect 14700 26460 14756 26516
rect 14588 26236 14644 26292
rect 15260 26290 15316 26292
rect 15260 26238 15262 26290
rect 15262 26238 15314 26290
rect 15314 26238 15316 26290
rect 15260 26236 15316 26238
rect 14700 25900 14756 25956
rect 14924 25618 14980 25620
rect 14924 25566 14926 25618
rect 14926 25566 14978 25618
rect 14978 25566 14980 25618
rect 14924 25564 14980 25566
rect 14812 25394 14868 25396
rect 14812 25342 14814 25394
rect 14814 25342 14866 25394
rect 14866 25342 14868 25394
rect 14812 25340 14868 25342
rect 15036 25394 15092 25396
rect 15036 25342 15038 25394
rect 15038 25342 15090 25394
rect 15090 25342 15092 25394
rect 15036 25340 15092 25342
rect 15260 25116 15316 25172
rect 14924 25004 14980 25060
rect 14588 23772 14644 23828
rect 14588 23548 14644 23604
rect 14812 24556 14868 24612
rect 14364 22482 14420 22484
rect 14364 22430 14366 22482
rect 14366 22430 14418 22482
rect 14418 22430 14420 22482
rect 14364 22428 14420 22430
rect 14140 21084 14196 21140
rect 14476 21532 14532 21588
rect 14364 20802 14420 20804
rect 14364 20750 14366 20802
rect 14366 20750 14418 20802
rect 14418 20750 14420 20802
rect 14364 20748 14420 20750
rect 14700 22092 14756 22148
rect 15260 23266 15316 23268
rect 15260 23214 15262 23266
rect 15262 23214 15314 23266
rect 15314 23214 15316 23266
rect 15260 23212 15316 23214
rect 15260 22764 15316 22820
rect 14588 20972 14644 21028
rect 14364 20412 14420 20468
rect 14028 19458 14084 19460
rect 14028 19406 14030 19458
rect 14030 19406 14082 19458
rect 14082 19406 14084 19458
rect 14028 19404 14084 19406
rect 13020 19292 13076 19348
rect 12124 19234 12180 19236
rect 12124 19182 12126 19234
rect 12126 19182 12178 19234
rect 12178 19182 12180 19234
rect 12124 19180 12180 19182
rect 12012 18508 12068 18564
rect 13804 19346 13860 19348
rect 13804 19294 13806 19346
rect 13806 19294 13858 19346
rect 13858 19294 13860 19346
rect 13804 19292 13860 19294
rect 13916 19180 13972 19236
rect 13804 17276 13860 17332
rect 11788 17164 11844 17220
rect 12908 16098 12964 16100
rect 12908 16046 12910 16098
rect 12910 16046 12962 16098
rect 12962 16046 12964 16098
rect 12908 16044 12964 16046
rect 13244 16044 13300 16100
rect 13132 15820 13188 15876
rect 11788 15260 11844 15316
rect 12460 15596 12516 15652
rect 12796 15538 12852 15540
rect 12796 15486 12798 15538
rect 12798 15486 12850 15538
rect 12850 15486 12852 15538
rect 12796 15484 12852 15486
rect 14028 16828 14084 16884
rect 14028 16156 14084 16212
rect 13468 15874 13524 15876
rect 13468 15822 13470 15874
rect 13470 15822 13522 15874
rect 13522 15822 13524 15874
rect 13468 15820 13524 15822
rect 12012 14642 12068 14644
rect 12012 14590 12014 14642
rect 12014 14590 12066 14642
rect 12066 14590 12068 14642
rect 12012 14588 12068 14590
rect 10780 14140 10836 14196
rect 11228 14140 11284 14196
rect 9436 11116 9492 11172
rect 8764 9826 8820 9828
rect 8764 9774 8766 9826
rect 8766 9774 8818 9826
rect 8818 9774 8820 9826
rect 8764 9772 8820 9774
rect 9772 11676 9828 11732
rect 9660 9772 9716 9828
rect 12460 14588 12516 14644
rect 10444 12908 10500 12964
rect 11452 12962 11508 12964
rect 11452 12910 11454 12962
rect 11454 12910 11506 12962
rect 11506 12910 11508 12962
rect 11452 12908 11508 12910
rect 11452 12236 11508 12292
rect 11676 12402 11732 12404
rect 11676 12350 11678 12402
rect 11678 12350 11730 12402
rect 11730 12350 11732 12402
rect 11676 12348 11732 12350
rect 11564 11564 11620 11620
rect 12124 12402 12180 12404
rect 12124 12350 12126 12402
rect 12126 12350 12178 12402
rect 12178 12350 12180 12402
rect 12124 12348 12180 12350
rect 13916 14306 13972 14308
rect 13916 14254 13918 14306
rect 13918 14254 13970 14306
rect 13970 14254 13972 14306
rect 13916 14252 13972 14254
rect 14588 20412 14644 20468
rect 15148 21756 15204 21812
rect 14924 21196 14980 21252
rect 15148 20412 15204 20468
rect 15484 25116 15540 25172
rect 15484 24780 15540 24836
rect 15932 28418 15988 28420
rect 15932 28366 15934 28418
rect 15934 28366 15986 28418
rect 15986 28366 15988 28418
rect 15932 28364 15988 28366
rect 16268 28700 16324 28756
rect 16380 28642 16436 28644
rect 16380 28590 16382 28642
rect 16382 28590 16434 28642
rect 16434 28590 16436 28642
rect 16380 28588 16436 28590
rect 16492 29260 16548 29316
rect 15820 27244 15876 27300
rect 15820 25788 15876 25844
rect 15932 25676 15988 25732
rect 16044 26348 16100 26404
rect 15932 25394 15988 25396
rect 15932 25342 15934 25394
rect 15934 25342 15986 25394
rect 15986 25342 15988 25394
rect 15932 25340 15988 25342
rect 16380 27970 16436 27972
rect 16380 27918 16382 27970
rect 16382 27918 16434 27970
rect 16434 27918 16436 27970
rect 16380 27916 16436 27918
rect 16380 26684 16436 26740
rect 16268 26402 16324 26404
rect 16268 26350 16270 26402
rect 16270 26350 16322 26402
rect 16322 26350 16324 26402
rect 16268 26348 16324 26350
rect 16716 29650 16772 29652
rect 16716 29598 16718 29650
rect 16718 29598 16770 29650
rect 16770 29598 16772 29650
rect 16716 29596 16772 29598
rect 16604 28364 16660 28420
rect 17052 28140 17108 28196
rect 16828 27916 16884 27972
rect 16716 27692 16772 27748
rect 16604 27132 16660 27188
rect 16940 26850 16996 26852
rect 16940 26798 16942 26850
rect 16942 26798 16994 26850
rect 16994 26798 16996 26850
rect 16940 26796 16996 26798
rect 16716 26460 16772 26516
rect 16156 24556 16212 24612
rect 17388 30828 17444 30884
rect 17388 29596 17444 29652
rect 17388 28418 17444 28420
rect 17388 28366 17390 28418
rect 17390 28366 17442 28418
rect 17442 28366 17444 28418
rect 17388 28364 17444 28366
rect 17276 26124 17332 26180
rect 17388 28140 17444 28196
rect 16716 25788 16772 25844
rect 16604 25676 16660 25732
rect 16492 25618 16548 25620
rect 16492 25566 16494 25618
rect 16494 25566 16546 25618
rect 16546 25566 16548 25618
rect 16492 25564 16548 25566
rect 16492 25004 16548 25060
rect 16940 25676 16996 25732
rect 16380 24556 16436 24612
rect 16716 24722 16772 24724
rect 16716 24670 16718 24722
rect 16718 24670 16770 24722
rect 16770 24670 16772 24722
rect 16716 24668 16772 24670
rect 16604 24444 16660 24500
rect 16492 23826 16548 23828
rect 16492 23774 16494 23826
rect 16494 23774 16546 23826
rect 16546 23774 16548 23826
rect 16492 23772 16548 23774
rect 16156 23212 16212 23268
rect 15820 22764 15876 22820
rect 16380 23100 16436 23156
rect 15708 22540 15764 22596
rect 15596 22428 15652 22484
rect 15372 21980 15428 22036
rect 15708 21756 15764 21812
rect 15596 21420 15652 21476
rect 15596 20860 15652 20916
rect 15372 20130 15428 20132
rect 15372 20078 15374 20130
rect 15374 20078 15426 20130
rect 15426 20078 15428 20130
rect 15372 20076 15428 20078
rect 15260 19292 15316 19348
rect 14812 18284 14868 18340
rect 14252 15820 14308 15876
rect 14700 15820 14756 15876
rect 15148 18674 15204 18676
rect 15148 18622 15150 18674
rect 15150 18622 15202 18674
rect 15202 18622 15204 18674
rect 15148 18620 15204 18622
rect 15036 16828 15092 16884
rect 14924 15484 14980 15540
rect 14588 15372 14644 15428
rect 14476 14924 14532 14980
rect 15372 15986 15428 15988
rect 15372 15934 15374 15986
rect 15374 15934 15426 15986
rect 15426 15934 15428 15986
rect 15372 15932 15428 15934
rect 15260 15596 15316 15652
rect 15260 14418 15316 14420
rect 15260 14366 15262 14418
rect 15262 14366 15314 14418
rect 15314 14366 15316 14418
rect 15260 14364 15316 14366
rect 14252 14306 14308 14308
rect 14252 14254 14254 14306
rect 14254 14254 14306 14306
rect 14306 14254 14308 14306
rect 14252 14252 14308 14254
rect 12684 12962 12740 12964
rect 12684 12910 12686 12962
rect 12686 12910 12738 12962
rect 12738 12910 12740 12962
rect 12684 12908 12740 12910
rect 13356 12290 13412 12292
rect 13356 12238 13358 12290
rect 13358 12238 13410 12290
rect 13410 12238 13412 12290
rect 13356 12236 13412 12238
rect 12796 11564 12852 11620
rect 14588 12962 14644 12964
rect 14588 12910 14590 12962
rect 14590 12910 14642 12962
rect 14642 12910 14644 12962
rect 14588 12908 14644 12910
rect 13916 12236 13972 12292
rect 11788 11116 11844 11172
rect 9884 9660 9940 9716
rect 11676 9884 11732 9940
rect 9660 9212 9716 9268
rect 12012 10332 12068 10388
rect 11788 9266 11844 9268
rect 11788 9214 11790 9266
rect 11790 9214 11842 9266
rect 11842 9214 11844 9266
rect 11788 9212 11844 9214
rect 12460 9996 12516 10052
rect 12124 9938 12180 9940
rect 12124 9886 12126 9938
rect 12126 9886 12178 9938
rect 12178 9886 12180 9938
rect 12124 9884 12180 9886
rect 8764 4060 8820 4116
rect 9772 4114 9828 4116
rect 9772 4062 9774 4114
rect 9774 4062 9826 4114
rect 9826 4062 9828 4114
rect 9772 4060 9828 4062
rect 12684 9212 12740 9268
rect 14140 9884 14196 9940
rect 15148 11676 15204 11732
rect 14812 11564 14868 11620
rect 15708 17276 15764 17332
rect 15596 15372 15652 15428
rect 15484 11676 15540 11732
rect 16044 21868 16100 21924
rect 16156 21196 16212 21252
rect 16716 22092 16772 22148
rect 16716 21756 16772 21812
rect 16268 20748 16324 20804
rect 16380 21308 16436 21364
rect 16156 20412 16212 20468
rect 15932 20188 15988 20244
rect 16604 21196 16660 21252
rect 16716 20188 16772 20244
rect 16380 19292 16436 19348
rect 16156 16604 16212 16660
rect 17612 32508 17668 32564
rect 17612 32338 17668 32340
rect 17612 32286 17614 32338
rect 17614 32286 17666 32338
rect 17666 32286 17668 32338
rect 17612 32284 17668 32286
rect 18284 34076 18340 34132
rect 18508 33964 18564 34020
rect 19292 35420 19348 35476
rect 19180 34690 19236 34692
rect 19180 34638 19182 34690
rect 19182 34638 19234 34690
rect 19234 34638 19236 34690
rect 19180 34636 19236 34638
rect 18508 33346 18564 33348
rect 18508 33294 18510 33346
rect 18510 33294 18562 33346
rect 18562 33294 18564 33346
rect 18508 33292 18564 33294
rect 18060 31724 18116 31780
rect 18508 31612 18564 31668
rect 18172 31106 18228 31108
rect 18172 31054 18174 31106
rect 18174 31054 18226 31106
rect 18226 31054 18228 31106
rect 18172 31052 18228 31054
rect 18060 30156 18116 30212
rect 17836 29932 17892 29988
rect 17612 29314 17668 29316
rect 17612 29262 17614 29314
rect 17614 29262 17666 29314
rect 17666 29262 17668 29314
rect 17612 29260 17668 29262
rect 17948 29260 18004 29316
rect 18508 29708 18564 29764
rect 18060 28588 18116 28644
rect 18172 28812 18228 28868
rect 17836 28252 17892 28308
rect 17500 27858 17556 27860
rect 17500 27806 17502 27858
rect 17502 27806 17554 27858
rect 17554 27806 17556 27858
rect 17500 27804 17556 27806
rect 17500 27244 17556 27300
rect 17948 27970 18004 27972
rect 17948 27918 17950 27970
rect 17950 27918 18002 27970
rect 18002 27918 18004 27970
rect 17948 27916 18004 27918
rect 17164 25004 17220 25060
rect 17276 24444 17332 24500
rect 17164 23660 17220 23716
rect 17388 23548 17444 23604
rect 17276 23324 17332 23380
rect 17612 26684 17668 26740
rect 17724 25900 17780 25956
rect 17612 25676 17668 25732
rect 17612 24946 17668 24948
rect 17612 24894 17614 24946
rect 17614 24894 17666 24946
rect 17666 24894 17668 24946
rect 17612 24892 17668 24894
rect 17500 23154 17556 23156
rect 17500 23102 17502 23154
rect 17502 23102 17554 23154
rect 17554 23102 17556 23154
rect 17500 23100 17556 23102
rect 17276 20524 17332 20580
rect 17724 23100 17780 23156
rect 17612 18338 17668 18340
rect 17612 18286 17614 18338
rect 17614 18286 17666 18338
rect 17666 18286 17668 18338
rect 17612 18284 17668 18286
rect 17052 16716 17108 16772
rect 17500 16828 17556 16884
rect 17388 16604 17444 16660
rect 16940 15932 16996 15988
rect 16156 14476 16212 14532
rect 16380 14476 16436 14532
rect 15932 14140 15988 14196
rect 17724 16156 17780 16212
rect 16492 14140 16548 14196
rect 17388 13020 17444 13076
rect 16716 12962 16772 12964
rect 16716 12910 16718 12962
rect 16718 12910 16770 12962
rect 16770 12910 16772 12962
rect 16716 12908 16772 12910
rect 15820 11564 15876 11620
rect 15596 11452 15652 11508
rect 16492 11506 16548 11508
rect 16492 11454 16494 11506
rect 16494 11454 16546 11506
rect 16546 11454 16548 11506
rect 16492 11452 16548 11454
rect 14364 9826 14420 9828
rect 14364 9774 14366 9826
rect 14366 9774 14418 9826
rect 14418 9774 14420 9826
rect 14364 9772 14420 9774
rect 15820 10780 15876 10836
rect 15372 10386 15428 10388
rect 15372 10334 15374 10386
rect 15374 10334 15426 10386
rect 15426 10334 15428 10386
rect 15372 10332 15428 10334
rect 15372 9938 15428 9940
rect 15372 9886 15374 9938
rect 15374 9886 15426 9938
rect 15426 9886 15428 9938
rect 15372 9884 15428 9886
rect 15708 9826 15764 9828
rect 15708 9774 15710 9826
rect 15710 9774 15762 9826
rect 15762 9774 15764 9826
rect 15708 9772 15764 9774
rect 14812 9212 14868 9268
rect 15932 9266 15988 9268
rect 15932 9214 15934 9266
rect 15934 9214 15986 9266
rect 15986 9214 15988 9266
rect 15932 9212 15988 9214
rect 12796 4060 12852 4116
rect 14028 4114 14084 4116
rect 14028 4062 14030 4114
rect 14030 4062 14082 4114
rect 14082 4062 14084 4114
rect 14028 4060 14084 4062
rect 16492 10834 16548 10836
rect 16492 10782 16494 10834
rect 16494 10782 16546 10834
rect 16546 10782 16548 10834
rect 16492 10780 16548 10782
rect 16940 9212 16996 9268
rect 17388 9660 17444 9716
rect 16828 6636 16884 6692
rect 17948 24892 18004 24948
rect 18508 28364 18564 28420
rect 18508 28028 18564 28084
rect 18284 27916 18340 27972
rect 18172 27074 18228 27076
rect 18172 27022 18174 27074
rect 18174 27022 18226 27074
rect 18226 27022 18228 27074
rect 18172 27020 18228 27022
rect 18396 27244 18452 27300
rect 18844 31052 18900 31108
rect 18956 33180 19012 33236
rect 20076 36988 20132 37044
rect 20300 36876 20356 36932
rect 19852 36258 19908 36260
rect 19852 36206 19854 36258
rect 19854 36206 19906 36258
rect 19906 36206 19908 36258
rect 19852 36204 19908 36206
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19740 35810 19796 35812
rect 19740 35758 19742 35810
rect 19742 35758 19794 35810
rect 19794 35758 19796 35810
rect 19740 35756 19796 35758
rect 21420 37212 21476 37268
rect 20860 36594 20916 36596
rect 20860 36542 20862 36594
rect 20862 36542 20914 36594
rect 20914 36542 20916 36594
rect 20860 36540 20916 36542
rect 21196 36316 21252 36372
rect 21868 43036 21924 43092
rect 22428 42252 22484 42308
rect 21756 42140 21812 42196
rect 22204 42140 22260 42196
rect 22652 42140 22708 42196
rect 25228 45890 25284 45892
rect 25228 45838 25230 45890
rect 25230 45838 25282 45890
rect 25282 45838 25284 45890
rect 25228 45836 25284 45838
rect 28252 46060 28308 46116
rect 29484 46114 29540 46116
rect 29484 46062 29486 46114
rect 29486 46062 29538 46114
rect 29538 46062 29540 46114
rect 29484 46060 29540 46062
rect 26908 45276 26964 45332
rect 28140 45330 28196 45332
rect 28140 45278 28142 45330
rect 28142 45278 28194 45330
rect 28194 45278 28196 45330
rect 28140 45276 28196 45278
rect 28476 45276 28532 45332
rect 25900 45218 25956 45220
rect 25900 45166 25902 45218
rect 25902 45166 25954 45218
rect 25954 45166 25956 45218
rect 25900 45164 25956 45166
rect 24220 44492 24276 44548
rect 24332 45052 24388 45108
rect 23996 43036 24052 43092
rect 25564 45106 25620 45108
rect 25564 45054 25566 45106
rect 25566 45054 25618 45106
rect 25618 45054 25620 45106
rect 25564 45052 25620 45054
rect 27132 45106 27188 45108
rect 27132 45054 27134 45106
rect 27134 45054 27186 45106
rect 27186 45054 27188 45106
rect 27132 45052 27188 45054
rect 25452 44546 25508 44548
rect 25452 44494 25454 44546
rect 25454 44494 25506 44546
rect 25506 44494 25508 44546
rect 25452 44492 25508 44494
rect 27468 44434 27524 44436
rect 27468 44382 27470 44434
rect 27470 44382 27522 44434
rect 27522 44382 27524 44434
rect 27468 44380 27524 44382
rect 27916 44434 27972 44436
rect 27916 44382 27918 44434
rect 27918 44382 27970 44434
rect 27970 44382 27972 44434
rect 27916 44380 27972 44382
rect 24444 44322 24500 44324
rect 24444 44270 24446 44322
rect 24446 44270 24498 44322
rect 24498 44270 24500 44322
rect 24444 44268 24500 44270
rect 24780 43036 24836 43092
rect 23884 42476 23940 42532
rect 22540 41074 22596 41076
rect 22540 41022 22542 41074
rect 22542 41022 22594 41074
rect 22594 41022 22596 41074
rect 22540 41020 22596 41022
rect 22316 40962 22372 40964
rect 22316 40910 22318 40962
rect 22318 40910 22370 40962
rect 22370 40910 22372 40962
rect 22316 40908 22372 40910
rect 22652 40962 22708 40964
rect 22652 40910 22654 40962
rect 22654 40910 22706 40962
rect 22706 40910 22708 40962
rect 22652 40908 22708 40910
rect 22876 41356 22932 41412
rect 23436 42140 23492 42196
rect 23548 41356 23604 41412
rect 22988 41244 23044 41300
rect 23884 41804 23940 41860
rect 26012 42140 26068 42196
rect 30940 46060 30996 46116
rect 29596 44492 29652 44548
rect 28252 43372 28308 43428
rect 28476 42754 28532 42756
rect 28476 42702 28478 42754
rect 28478 42702 28530 42754
rect 28530 42702 28532 42754
rect 28476 42700 28532 42702
rect 29036 43426 29092 43428
rect 29036 43374 29038 43426
rect 29038 43374 29090 43426
rect 29090 43374 29092 43426
rect 29036 43372 29092 43374
rect 28140 42028 28196 42084
rect 28924 42924 28980 42980
rect 25340 41916 25396 41972
rect 23772 41298 23828 41300
rect 23772 41246 23774 41298
rect 23774 41246 23826 41298
rect 23826 41246 23828 41298
rect 23772 41244 23828 41246
rect 23100 41074 23156 41076
rect 23100 41022 23102 41074
rect 23102 41022 23154 41074
rect 23154 41022 23156 41074
rect 23100 41020 23156 41022
rect 22092 40572 22148 40628
rect 21980 39506 22036 39508
rect 21980 39454 21982 39506
rect 21982 39454 22034 39506
rect 22034 39454 22036 39506
rect 21980 39452 22036 39454
rect 21644 39394 21700 39396
rect 21644 39342 21646 39394
rect 21646 39342 21698 39394
rect 21698 39342 21700 39394
rect 21644 39340 21700 39342
rect 21756 37772 21812 37828
rect 22316 39564 22372 39620
rect 22428 39340 22484 39396
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19964 34018 20020 34020
rect 19964 33966 19966 34018
rect 19966 33966 20018 34018
rect 20018 33966 20020 34018
rect 19964 33964 20020 33966
rect 19628 32956 19684 33012
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19404 31890 19460 31892
rect 19404 31838 19406 31890
rect 19406 31838 19458 31890
rect 19458 31838 19460 31890
rect 19404 31836 19460 31838
rect 19068 31724 19124 31780
rect 19068 31554 19124 31556
rect 19068 31502 19070 31554
rect 19070 31502 19122 31554
rect 19122 31502 19124 31554
rect 19068 31500 19124 31502
rect 19516 31164 19572 31220
rect 19404 31052 19460 31108
rect 18956 30044 19012 30100
rect 19180 30268 19236 30324
rect 18956 29820 19012 29876
rect 18956 29314 19012 29316
rect 18956 29262 18958 29314
rect 18958 29262 19010 29314
rect 19010 29262 19012 29314
rect 18956 29260 19012 29262
rect 19180 29986 19236 29988
rect 19180 29934 19182 29986
rect 19182 29934 19234 29986
rect 19234 29934 19236 29986
rect 19180 29932 19236 29934
rect 18620 26908 18676 26964
rect 18732 28924 18788 28980
rect 18508 26684 18564 26740
rect 17948 23324 18004 23380
rect 18172 26124 18228 26180
rect 18956 28588 19012 28644
rect 18844 28252 18900 28308
rect 19852 31836 19908 31892
rect 19740 31778 19796 31780
rect 19740 31726 19742 31778
rect 19742 31726 19794 31778
rect 19794 31726 19796 31778
rect 19740 31724 19796 31726
rect 19964 31778 20020 31780
rect 19964 31726 19966 31778
rect 19966 31726 20018 31778
rect 20018 31726 20020 31778
rect 19964 31724 20020 31726
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20300 31276 20356 31332
rect 20412 31164 20468 31220
rect 20300 31106 20356 31108
rect 20300 31054 20302 31106
rect 20302 31054 20354 31106
rect 20354 31054 20356 31106
rect 20300 31052 20356 31054
rect 19516 30380 19572 30436
rect 19628 30604 19684 30660
rect 19404 29708 19460 29764
rect 19740 30322 19796 30324
rect 19740 30270 19742 30322
rect 19742 30270 19794 30322
rect 19794 30270 19796 30322
rect 19740 30268 19796 30270
rect 20636 30994 20692 30996
rect 20636 30942 20638 30994
rect 20638 30942 20690 30994
rect 20690 30942 20692 30994
rect 20636 30940 20692 30942
rect 20524 30380 20580 30436
rect 20412 30268 20468 30324
rect 20188 30044 20244 30100
rect 20076 29986 20132 29988
rect 20076 29934 20078 29986
rect 20078 29934 20130 29986
rect 20130 29934 20132 29986
rect 20076 29932 20132 29934
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19628 29426 19684 29428
rect 19628 29374 19630 29426
rect 19630 29374 19682 29426
rect 19682 29374 19684 29426
rect 19628 29372 19684 29374
rect 19516 29260 19572 29316
rect 20636 30044 20692 30100
rect 20412 29314 20468 29316
rect 20412 29262 20414 29314
rect 20414 29262 20466 29314
rect 20466 29262 20468 29314
rect 20412 29260 20468 29262
rect 21084 29260 21140 29316
rect 19292 28924 19348 28980
rect 19404 29148 19460 29204
rect 19180 26796 19236 26852
rect 19292 28364 19348 28420
rect 19292 27132 19348 27188
rect 18956 26236 19012 26292
rect 18620 25340 18676 25396
rect 18396 25282 18452 25284
rect 18396 25230 18398 25282
rect 18398 25230 18450 25282
rect 18450 25230 18452 25282
rect 18396 25228 18452 25230
rect 18508 25116 18564 25172
rect 18284 24556 18340 24612
rect 18620 24722 18676 24724
rect 18620 24670 18622 24722
rect 18622 24670 18674 24722
rect 18674 24670 18676 24722
rect 18620 24668 18676 24670
rect 18508 24556 18564 24612
rect 18172 23324 18228 23380
rect 17948 23100 18004 23156
rect 17948 22204 18004 22260
rect 18060 22092 18116 22148
rect 18060 19964 18116 20020
rect 18284 22092 18340 22148
rect 18844 24780 18900 24836
rect 19068 25004 19124 25060
rect 18732 22428 18788 22484
rect 18844 23324 18900 23380
rect 18396 21420 18452 21476
rect 18172 18562 18228 18564
rect 18172 18510 18174 18562
rect 18174 18510 18226 18562
rect 18226 18510 18228 18562
rect 18172 18508 18228 18510
rect 18620 18508 18676 18564
rect 17948 18284 18004 18340
rect 18060 18226 18116 18228
rect 18060 18174 18062 18226
rect 18062 18174 18114 18226
rect 18114 18174 18116 18226
rect 18060 18172 18116 18174
rect 18396 17724 18452 17780
rect 19404 27244 19460 27300
rect 19628 29148 19684 29204
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19852 27970 19908 27972
rect 19852 27918 19854 27970
rect 19854 27918 19906 27970
rect 19906 27918 19908 27970
rect 19852 27916 19908 27918
rect 20412 27970 20468 27972
rect 20412 27918 20414 27970
rect 20414 27918 20466 27970
rect 20466 27918 20468 27970
rect 20412 27916 20468 27918
rect 20524 27804 20580 27860
rect 19964 27692 20020 27748
rect 19964 27244 20020 27300
rect 20524 27244 20580 27300
rect 20412 27074 20468 27076
rect 20412 27022 20414 27074
rect 20414 27022 20466 27074
rect 20466 27022 20468 27074
rect 20412 27020 20468 27022
rect 20300 26796 20356 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19852 26236 19908 26292
rect 19964 26460 20020 26516
rect 20300 26460 20356 26516
rect 20188 26124 20244 26180
rect 19740 25228 19796 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19180 24610 19236 24612
rect 19180 24558 19182 24610
rect 19182 24558 19234 24610
rect 19234 24558 19236 24610
rect 19180 24556 19236 24558
rect 19180 23772 19236 23828
rect 19068 21756 19124 21812
rect 19852 24834 19908 24836
rect 19852 24782 19854 24834
rect 19854 24782 19906 24834
rect 19906 24782 19908 24834
rect 19852 24780 19908 24782
rect 20412 24892 20468 24948
rect 20188 23772 20244 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19404 22428 19460 22484
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19852 21698 19908 21700
rect 19852 21646 19854 21698
rect 19854 21646 19906 21698
rect 19906 21646 19908 21698
rect 19852 21644 19908 21646
rect 19404 21586 19460 21588
rect 19404 21534 19406 21586
rect 19406 21534 19458 21586
rect 19458 21534 19460 21586
rect 19404 21532 19460 21534
rect 19964 20636 20020 20692
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19404 18284 19460 18340
rect 19516 18172 19572 18228
rect 18844 17052 18900 17108
rect 19068 17500 19124 17556
rect 18508 16828 18564 16884
rect 17948 16210 18004 16212
rect 17948 16158 17950 16210
rect 17950 16158 18002 16210
rect 18002 16158 18004 16210
rect 17948 16156 18004 16158
rect 19404 17106 19460 17108
rect 19404 17054 19406 17106
rect 19406 17054 19458 17106
rect 19458 17054 19460 17106
rect 19404 17052 19460 17054
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19740 17500 19796 17556
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19852 17106 19908 17108
rect 19852 17054 19854 17106
rect 19854 17054 19906 17106
rect 19906 17054 19908 17106
rect 19852 17052 19908 17054
rect 19068 16716 19124 16772
rect 19068 16156 19124 16212
rect 20076 16994 20132 16996
rect 20076 16942 20078 16994
rect 20078 16942 20130 16994
rect 20130 16942 20132 16994
rect 20076 16940 20132 16942
rect 20300 22988 20356 23044
rect 20524 21474 20580 21476
rect 20524 21422 20526 21474
rect 20526 21422 20578 21474
rect 20578 21422 20580 21474
rect 20524 21420 20580 21422
rect 20748 25452 20804 25508
rect 20860 24892 20916 24948
rect 20860 23324 20916 23380
rect 22316 36370 22372 36372
rect 22316 36318 22318 36370
rect 22318 36318 22370 36370
rect 22370 36318 22372 36370
rect 22316 36316 22372 36318
rect 22204 35868 22260 35924
rect 21980 35532 22036 35588
rect 21644 34860 21700 34916
rect 21756 31836 21812 31892
rect 21532 31164 21588 31220
rect 21644 30492 21700 30548
rect 21756 28364 21812 28420
rect 21308 27468 21364 27524
rect 21308 27298 21364 27300
rect 21308 27246 21310 27298
rect 21310 27246 21362 27298
rect 21362 27246 21364 27298
rect 21308 27244 21364 27246
rect 21196 27020 21252 27076
rect 21196 26124 21252 26180
rect 22764 39452 22820 39508
rect 22652 36540 22708 36596
rect 22540 36258 22596 36260
rect 22540 36206 22542 36258
rect 22542 36206 22594 36258
rect 22594 36206 22596 36258
rect 22540 36204 22596 36206
rect 22876 35868 22932 35924
rect 22428 34914 22484 34916
rect 22428 34862 22430 34914
rect 22430 34862 22482 34914
rect 22482 34862 22484 34914
rect 22428 34860 22484 34862
rect 22316 34748 22372 34804
rect 21980 33628 22036 33684
rect 22316 28364 22372 28420
rect 21644 27020 21700 27076
rect 21980 27074 22036 27076
rect 21980 27022 21982 27074
rect 21982 27022 22034 27074
rect 22034 27022 22036 27074
rect 21980 27020 22036 27022
rect 21532 26460 21588 26516
rect 21420 26236 21476 26292
rect 21756 26572 21812 26628
rect 21980 26796 22036 26852
rect 21980 26290 22036 26292
rect 21980 26238 21982 26290
rect 21982 26238 22034 26290
rect 22034 26238 22036 26290
rect 21980 26236 22036 26238
rect 21868 25900 21924 25956
rect 22092 26012 22148 26068
rect 21308 23436 21364 23492
rect 21084 22988 21140 23044
rect 20860 22146 20916 22148
rect 20860 22094 20862 22146
rect 20862 22094 20914 22146
rect 20914 22094 20916 22146
rect 20860 22092 20916 22094
rect 21308 22146 21364 22148
rect 21308 22094 21310 22146
rect 21310 22094 21362 22146
rect 21362 22094 21364 22146
rect 21308 22092 21364 22094
rect 20748 21868 20804 21924
rect 20748 21698 20804 21700
rect 20748 21646 20750 21698
rect 20750 21646 20802 21698
rect 20802 21646 20804 21698
rect 20748 21644 20804 21646
rect 21084 21420 21140 21476
rect 20412 20690 20468 20692
rect 20412 20638 20414 20690
rect 20414 20638 20466 20690
rect 20466 20638 20468 20690
rect 20412 20636 20468 20638
rect 20412 19628 20468 19684
rect 20300 17554 20356 17556
rect 20300 17502 20302 17554
rect 20302 17502 20354 17554
rect 20354 17502 20356 17554
rect 20300 17500 20356 17502
rect 20188 16268 20244 16324
rect 18956 15932 19012 15988
rect 19740 15932 19796 15988
rect 20076 16210 20132 16212
rect 20076 16158 20078 16210
rect 20078 16158 20130 16210
rect 20130 16158 20132 16210
rect 20076 16156 20132 16158
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19964 15260 20020 15316
rect 19404 15202 19460 15204
rect 19404 15150 19406 15202
rect 19406 15150 19458 15202
rect 19458 15150 19460 15202
rect 19404 15148 19460 15150
rect 19852 14700 19908 14756
rect 20076 15148 20132 15204
rect 21084 20300 21140 20356
rect 20748 19628 20804 19684
rect 20748 17778 20804 17780
rect 20748 17726 20750 17778
rect 20750 17726 20802 17778
rect 20802 17726 20804 17778
rect 20748 17724 20804 17726
rect 20860 17164 20916 17220
rect 20748 16994 20804 16996
rect 20748 16942 20750 16994
rect 20750 16942 20802 16994
rect 20802 16942 20804 16994
rect 20748 16940 20804 16942
rect 19068 14476 19124 14532
rect 18060 12012 18116 12068
rect 20076 14364 20132 14420
rect 19964 14306 20020 14308
rect 19964 14254 19966 14306
rect 19966 14254 20018 14306
rect 20018 14254 20020 14306
rect 19964 14252 20020 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20412 14364 20468 14420
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19180 12066 19236 12068
rect 19180 12014 19182 12066
rect 19182 12014 19234 12066
rect 19234 12014 19236 12066
rect 19180 12012 19236 12014
rect 20524 13692 20580 13748
rect 20300 13580 20356 13636
rect 20300 13074 20356 13076
rect 20300 13022 20302 13074
rect 20302 13022 20354 13074
rect 20354 13022 20356 13074
rect 20300 13020 20356 13022
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20524 12290 20580 12292
rect 20524 12238 20526 12290
rect 20526 12238 20578 12290
rect 20578 12238 20580 12290
rect 20524 12236 20580 12238
rect 19404 10722 19460 10724
rect 19404 10670 19406 10722
rect 19406 10670 19458 10722
rect 19458 10670 19460 10722
rect 19404 10668 19460 10670
rect 20076 10668 20132 10724
rect 18620 9660 18676 9716
rect 21308 20018 21364 20020
rect 21308 19966 21310 20018
rect 21310 19966 21362 20018
rect 21362 19966 21364 20018
rect 21308 19964 21364 19966
rect 21532 23212 21588 23268
rect 21868 23212 21924 23268
rect 21644 21586 21700 21588
rect 21644 21534 21646 21586
rect 21646 21534 21698 21586
rect 21698 21534 21700 21586
rect 21644 21532 21700 21534
rect 21980 20300 22036 20356
rect 21532 19068 21588 19124
rect 21420 18338 21476 18340
rect 21420 18286 21422 18338
rect 21422 18286 21474 18338
rect 21474 18286 21476 18338
rect 21420 18284 21476 18286
rect 21532 17724 21588 17780
rect 21308 17612 21364 17668
rect 21308 16268 21364 16324
rect 20972 15314 21028 15316
rect 20972 15262 20974 15314
rect 20974 15262 21026 15314
rect 21026 15262 21028 15314
rect 20972 15260 21028 15262
rect 21196 14812 21252 14868
rect 20972 14252 21028 14308
rect 20860 13746 20916 13748
rect 20860 13694 20862 13746
rect 20862 13694 20914 13746
rect 20914 13694 20916 13746
rect 20860 13692 20916 13694
rect 20972 12012 21028 12068
rect 20748 11394 20804 11396
rect 20748 11342 20750 11394
rect 20750 11342 20802 11394
rect 20802 11342 20804 11394
rect 20748 11340 20804 11342
rect 21420 15932 21476 15988
rect 21420 15314 21476 15316
rect 21420 15262 21422 15314
rect 21422 15262 21474 15314
rect 21474 15262 21476 15314
rect 21420 15260 21476 15262
rect 21420 14306 21476 14308
rect 21420 14254 21422 14306
rect 21422 14254 21474 14306
rect 21474 14254 21476 14306
rect 21420 14252 21476 14254
rect 21644 17612 21700 17668
rect 22876 34914 22932 34916
rect 22876 34862 22878 34914
rect 22878 34862 22930 34914
rect 22930 34862 22932 34914
rect 22876 34860 22932 34862
rect 23212 39564 23268 39620
rect 23772 39506 23828 39508
rect 23772 39454 23774 39506
rect 23774 39454 23826 39506
rect 23826 39454 23828 39506
rect 23772 39452 23828 39454
rect 23996 38892 24052 38948
rect 25228 40908 25284 40964
rect 25004 40348 25060 40404
rect 24668 38834 24724 38836
rect 24668 38782 24670 38834
rect 24670 38782 24722 38834
rect 24722 38782 24724 38834
rect 24668 38780 24724 38782
rect 23212 37772 23268 37828
rect 23548 36988 23604 37044
rect 23548 35644 23604 35700
rect 23324 35586 23380 35588
rect 23324 35534 23326 35586
rect 23326 35534 23378 35586
rect 23378 35534 23380 35586
rect 23324 35532 23380 35534
rect 23212 34748 23268 34804
rect 23324 34636 23380 34692
rect 23100 33628 23156 33684
rect 22876 33404 22932 33460
rect 22652 33180 22708 33236
rect 22988 33234 23044 33236
rect 22988 33182 22990 33234
rect 22990 33182 23042 33234
rect 23042 33182 23044 33234
rect 22988 33180 23044 33182
rect 23212 31836 23268 31892
rect 22764 31276 22820 31332
rect 23212 31218 23268 31220
rect 23212 31166 23214 31218
rect 23214 31166 23266 31218
rect 23266 31166 23268 31218
rect 23212 31164 23268 31166
rect 22652 30492 22708 30548
rect 24892 35138 24948 35140
rect 24892 35086 24894 35138
rect 24894 35086 24946 35138
rect 24946 35086 24948 35138
rect 24892 35084 24948 35086
rect 24556 34748 24612 34804
rect 24444 34300 24500 34356
rect 25004 34076 25060 34132
rect 24332 33628 24388 33684
rect 27916 41970 27972 41972
rect 27916 41918 27918 41970
rect 27918 41918 27970 41970
rect 27970 41918 27972 41970
rect 27916 41916 27972 41918
rect 27580 41804 27636 41860
rect 25340 38780 25396 38836
rect 26124 41132 26180 41188
rect 27580 41186 27636 41188
rect 27580 41134 27582 41186
rect 27582 41134 27634 41186
rect 27634 41134 27636 41186
rect 27580 41132 27636 41134
rect 27132 40908 27188 40964
rect 26572 40684 26628 40740
rect 27020 40514 27076 40516
rect 27020 40462 27022 40514
rect 27022 40462 27074 40514
rect 27074 40462 27076 40514
rect 27020 40460 27076 40462
rect 26908 40236 26964 40292
rect 27580 40684 27636 40740
rect 27132 39788 27188 39844
rect 26908 39564 26964 39620
rect 27580 40348 27636 40404
rect 27468 39788 27524 39844
rect 28476 41916 28532 41972
rect 28140 40908 28196 40964
rect 28476 41132 28532 41188
rect 28028 40236 28084 40292
rect 27916 39788 27972 39844
rect 28140 39730 28196 39732
rect 28140 39678 28142 39730
rect 28142 39678 28194 39730
rect 28194 39678 28196 39730
rect 28140 39676 28196 39678
rect 26460 39340 26516 39396
rect 26572 38722 26628 38724
rect 26572 38670 26574 38722
rect 26574 38670 26626 38722
rect 26626 38670 26628 38722
rect 26572 38668 26628 38670
rect 25340 34354 25396 34356
rect 25340 34302 25342 34354
rect 25342 34302 25394 34354
rect 25394 34302 25396 34354
rect 25340 34300 25396 34302
rect 25228 33404 25284 33460
rect 23660 31948 23716 32004
rect 23660 31500 23716 31556
rect 24108 30380 24164 30436
rect 22316 27298 22372 27300
rect 22316 27246 22318 27298
rect 22318 27246 22370 27298
rect 22370 27246 22372 27298
rect 22316 27244 22372 27246
rect 23100 27244 23156 27300
rect 22316 27074 22372 27076
rect 22316 27022 22318 27074
rect 22318 27022 22370 27074
rect 22370 27022 22372 27074
rect 22316 27020 22372 27022
rect 22540 26514 22596 26516
rect 22540 26462 22542 26514
rect 22542 26462 22594 26514
rect 22594 26462 22596 26514
rect 22540 26460 22596 26462
rect 22316 25340 22372 25396
rect 22204 23212 22260 23268
rect 22428 22652 22484 22708
rect 22204 22092 22260 22148
rect 22204 21810 22260 21812
rect 22204 21758 22206 21810
rect 22206 21758 22258 21810
rect 22258 21758 22260 21810
rect 22204 21756 22260 21758
rect 21980 17388 22036 17444
rect 21868 16882 21924 16884
rect 21868 16830 21870 16882
rect 21870 16830 21922 16882
rect 21922 16830 21924 16882
rect 21868 16828 21924 16830
rect 22316 20300 22372 20356
rect 22204 16604 22260 16660
rect 21644 16380 21700 16436
rect 21980 15932 22036 15988
rect 21644 15426 21700 15428
rect 21644 15374 21646 15426
rect 21646 15374 21698 15426
rect 21698 15374 21700 15426
rect 21644 15372 21700 15374
rect 22092 15426 22148 15428
rect 22092 15374 22094 15426
rect 22094 15374 22146 15426
rect 22146 15374 22148 15426
rect 22092 15372 22148 15374
rect 22316 15314 22372 15316
rect 22316 15262 22318 15314
rect 22318 15262 22370 15314
rect 22370 15262 22372 15314
rect 22316 15260 22372 15262
rect 22092 14924 22148 14980
rect 21644 14700 21700 14756
rect 21868 14530 21924 14532
rect 21868 14478 21870 14530
rect 21870 14478 21922 14530
rect 21922 14478 21924 14530
rect 21868 14476 21924 14478
rect 21532 13916 21588 13972
rect 21532 13634 21588 13636
rect 21532 13582 21534 13634
rect 21534 13582 21586 13634
rect 21586 13582 21588 13634
rect 21532 13580 21588 13582
rect 21756 13580 21812 13636
rect 21532 12962 21588 12964
rect 21532 12910 21534 12962
rect 21534 12910 21586 12962
rect 21586 12910 21588 12962
rect 21532 12908 21588 12910
rect 21756 13356 21812 13412
rect 21420 12236 21476 12292
rect 20076 9772 20132 9828
rect 20524 9772 20580 9828
rect 20188 9660 20244 9716
rect 20076 9602 20132 9604
rect 20076 9550 20078 9602
rect 20078 9550 20130 9602
rect 20130 9550 20132 9602
rect 20076 9548 20132 9550
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19740 9042 19796 9044
rect 19740 8990 19742 9042
rect 19742 8990 19794 9042
rect 19794 8990 19796 9042
rect 19740 8988 19796 8990
rect 19180 8876 19236 8932
rect 20076 8876 20132 8932
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20748 9154 20804 9156
rect 20748 9102 20750 9154
rect 20750 9102 20802 9154
rect 20802 9102 20804 9154
rect 20748 9100 20804 9102
rect 20524 8988 20580 9044
rect 21868 11340 21924 11396
rect 22540 21586 22596 21588
rect 22540 21534 22542 21586
rect 22542 21534 22594 21586
rect 22594 21534 22596 21586
rect 22540 21532 22596 21534
rect 22540 20802 22596 20804
rect 22540 20750 22542 20802
rect 22542 20750 22594 20802
rect 22594 20750 22596 20802
rect 22540 20748 22596 20750
rect 22988 26796 23044 26852
rect 22876 26572 22932 26628
rect 23100 26012 23156 26068
rect 22876 24780 22932 24836
rect 23436 27634 23492 27636
rect 23436 27582 23438 27634
rect 23438 27582 23490 27634
rect 23490 27582 23492 27634
rect 23436 27580 23492 27582
rect 23436 27132 23492 27188
rect 23324 27074 23380 27076
rect 23324 27022 23326 27074
rect 23326 27022 23378 27074
rect 23378 27022 23380 27074
rect 23324 27020 23380 27022
rect 23996 27580 24052 27636
rect 24108 27356 24164 27412
rect 23772 26796 23828 26852
rect 23884 27132 23940 27188
rect 23884 26908 23940 26964
rect 23436 26066 23492 26068
rect 23436 26014 23438 26066
rect 23438 26014 23490 26066
rect 23490 26014 23492 26066
rect 23436 26012 23492 26014
rect 22652 19964 22708 20020
rect 22764 23660 22820 23716
rect 22540 16994 22596 16996
rect 22540 16942 22542 16994
rect 22542 16942 22594 16994
rect 22594 16942 22596 16994
rect 22540 16940 22596 16942
rect 22652 15314 22708 15316
rect 22652 15262 22654 15314
rect 22654 15262 22706 15314
rect 22706 15262 22708 15314
rect 22652 15260 22708 15262
rect 22540 14252 22596 14308
rect 22428 9996 22484 10052
rect 21868 9826 21924 9828
rect 21868 9774 21870 9826
rect 21870 9774 21922 9826
rect 21922 9774 21924 9826
rect 21868 9772 21924 9774
rect 22204 9826 22260 9828
rect 22204 9774 22206 9826
rect 22206 9774 22258 9826
rect 22258 9774 22260 9826
rect 22204 9772 22260 9774
rect 23100 22146 23156 22148
rect 23100 22094 23102 22146
rect 23102 22094 23154 22146
rect 23154 22094 23156 22146
rect 23100 22092 23156 22094
rect 23436 25676 23492 25732
rect 23324 23826 23380 23828
rect 23324 23774 23326 23826
rect 23326 23774 23378 23826
rect 23378 23774 23380 23826
rect 23324 23772 23380 23774
rect 22876 21698 22932 21700
rect 22876 21646 22878 21698
rect 22878 21646 22930 21698
rect 22930 21646 22932 21698
rect 22876 21644 22932 21646
rect 23324 23436 23380 23492
rect 22988 21532 23044 21588
rect 22876 19628 22932 19684
rect 23212 21586 23268 21588
rect 23212 21534 23214 21586
rect 23214 21534 23266 21586
rect 23266 21534 23268 21586
rect 23212 21532 23268 21534
rect 23436 21308 23492 21364
rect 23324 20748 23380 20804
rect 24108 27074 24164 27076
rect 24108 27022 24110 27074
rect 24110 27022 24162 27074
rect 24162 27022 24164 27074
rect 24108 27020 24164 27022
rect 24444 32060 24500 32116
rect 25564 31612 25620 31668
rect 24444 30380 24500 30436
rect 25228 30434 25284 30436
rect 25228 30382 25230 30434
rect 25230 30382 25282 30434
rect 25282 30382 25284 30434
rect 25228 30380 25284 30382
rect 24556 30210 24612 30212
rect 24556 30158 24558 30210
rect 24558 30158 24610 30210
rect 24610 30158 24612 30210
rect 24556 30156 24612 30158
rect 24108 26796 24164 26852
rect 24332 26460 24388 26516
rect 23660 25788 23716 25844
rect 24108 26012 24164 26068
rect 23996 24834 24052 24836
rect 23996 24782 23998 24834
rect 23998 24782 24050 24834
rect 24050 24782 24052 24834
rect 23996 24780 24052 24782
rect 23996 24220 24052 24276
rect 23772 23826 23828 23828
rect 23772 23774 23774 23826
rect 23774 23774 23826 23826
rect 23826 23774 23828 23826
rect 23772 23772 23828 23774
rect 23772 22652 23828 22708
rect 23660 22092 23716 22148
rect 23660 21586 23716 21588
rect 23660 21534 23662 21586
rect 23662 21534 23714 21586
rect 23714 21534 23716 21586
rect 23660 21532 23716 21534
rect 23884 20860 23940 20916
rect 23100 17724 23156 17780
rect 23324 16380 23380 16436
rect 23772 19964 23828 20020
rect 24332 21532 24388 21588
rect 24220 20860 24276 20916
rect 24556 24220 24612 24276
rect 24668 29932 24724 29988
rect 24668 23772 24724 23828
rect 24892 26908 24948 26964
rect 25228 27074 25284 27076
rect 25228 27022 25230 27074
rect 25230 27022 25282 27074
rect 25282 27022 25284 27074
rect 25228 27020 25284 27022
rect 25004 26460 25060 26516
rect 25340 26796 25396 26852
rect 25676 26908 25732 26964
rect 25452 26348 25508 26404
rect 25340 25900 25396 25956
rect 25228 25788 25284 25844
rect 26908 39340 26964 39396
rect 27356 39228 27412 39284
rect 27020 38668 27076 38724
rect 26796 38444 26852 38500
rect 27356 39004 27412 39060
rect 27580 39116 27636 39172
rect 28588 40962 28644 40964
rect 28588 40910 28590 40962
rect 28590 40910 28642 40962
rect 28642 40910 28644 40962
rect 28588 40908 28644 40910
rect 28252 39004 28308 39060
rect 28588 40348 28644 40404
rect 28812 39788 28868 39844
rect 28812 39228 28868 39284
rect 28700 39058 28756 39060
rect 28700 39006 28702 39058
rect 28702 39006 28754 39058
rect 28754 39006 28756 39058
rect 28700 39004 28756 39006
rect 27132 37996 27188 38052
rect 27356 38556 27412 38612
rect 27244 36876 27300 36932
rect 26124 34242 26180 34244
rect 26124 34190 26126 34242
rect 26126 34190 26178 34242
rect 26178 34190 26180 34242
rect 26124 34188 26180 34190
rect 26796 34076 26852 34132
rect 26124 33964 26180 34020
rect 26012 30210 26068 30212
rect 26012 30158 26014 30210
rect 26014 30158 26066 30210
rect 26066 30158 26068 30210
rect 26012 30156 26068 30158
rect 25900 27020 25956 27076
rect 24668 23436 24724 23492
rect 24668 22092 24724 22148
rect 24668 21810 24724 21812
rect 24668 21758 24670 21810
rect 24670 21758 24722 21810
rect 24722 21758 24724 21810
rect 24668 21756 24724 21758
rect 24780 21420 24836 21476
rect 24556 20914 24612 20916
rect 24556 20862 24558 20914
rect 24558 20862 24610 20914
rect 24610 20862 24612 20914
rect 24556 20860 24612 20862
rect 25228 23436 25284 23492
rect 25228 21868 25284 21924
rect 25116 21532 25172 21588
rect 25340 21644 25396 21700
rect 25004 20748 25060 20804
rect 25340 21474 25396 21476
rect 25340 21422 25342 21474
rect 25342 21422 25394 21474
rect 25394 21422 25396 21474
rect 25340 21420 25396 21422
rect 25004 20578 25060 20580
rect 25004 20526 25006 20578
rect 25006 20526 25058 20578
rect 25058 20526 25060 20578
rect 25004 20524 25060 20526
rect 25564 23772 25620 23828
rect 25564 22146 25620 22148
rect 25564 22094 25566 22146
rect 25566 22094 25618 22146
rect 25618 22094 25620 22146
rect 25564 22092 25620 22094
rect 24668 20130 24724 20132
rect 24668 20078 24670 20130
rect 24670 20078 24722 20130
rect 24722 20078 24724 20130
rect 24668 20076 24724 20078
rect 25564 20914 25620 20916
rect 25564 20862 25566 20914
rect 25566 20862 25618 20914
rect 25618 20862 25620 20914
rect 25564 20860 25620 20862
rect 24556 19740 24612 19796
rect 23548 13580 23604 13636
rect 25452 20076 25508 20132
rect 25676 19068 25732 19124
rect 23548 11788 23604 11844
rect 23660 12684 23716 12740
rect 24556 17948 24612 18004
rect 25340 18060 25396 18116
rect 25676 17612 25732 17668
rect 25004 17164 25060 17220
rect 24668 17052 24724 17108
rect 24220 14812 24276 14868
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 23772 12012 23828 12068
rect 23660 11452 23716 11508
rect 25452 16882 25508 16884
rect 25452 16830 25454 16882
rect 25454 16830 25506 16882
rect 25506 16830 25508 16882
rect 25452 16828 25508 16830
rect 25228 16492 25284 16548
rect 25228 15596 25284 15652
rect 26236 33404 26292 33460
rect 26908 34076 26964 34132
rect 27916 38834 27972 38836
rect 27916 38782 27918 38834
rect 27918 38782 27970 38834
rect 27970 38782 27972 38834
rect 27916 38780 27972 38782
rect 28252 38668 28308 38724
rect 27692 38444 27748 38500
rect 27916 38556 27972 38612
rect 27916 37436 27972 37492
rect 28140 36876 28196 36932
rect 27020 33458 27076 33460
rect 27020 33406 27022 33458
rect 27022 33406 27074 33458
rect 27074 33406 27076 33458
rect 27020 33404 27076 33406
rect 26908 32844 26964 32900
rect 26796 32732 26852 32788
rect 26908 32620 26964 32676
rect 27580 33404 27636 33460
rect 28028 33404 28084 33460
rect 27692 33346 27748 33348
rect 27692 33294 27694 33346
rect 27694 33294 27746 33346
rect 27746 33294 27748 33346
rect 27692 33292 27748 33294
rect 27020 32396 27076 32452
rect 26908 31388 26964 31444
rect 26684 29260 26740 29316
rect 26236 28364 26292 28420
rect 26460 28588 26516 28644
rect 26236 27244 26292 27300
rect 26348 27186 26404 27188
rect 26348 27134 26350 27186
rect 26350 27134 26402 27186
rect 26402 27134 26404 27186
rect 26348 27132 26404 27134
rect 26572 26796 26628 26852
rect 26684 28364 26740 28420
rect 26124 21868 26180 21924
rect 26348 24780 26404 24836
rect 25900 21644 25956 21700
rect 26236 20748 26292 20804
rect 25900 19852 25956 19908
rect 26124 18060 26180 18116
rect 26012 17388 26068 17444
rect 26012 15596 26068 15652
rect 26908 28588 26964 28644
rect 26908 27298 26964 27300
rect 26908 27246 26910 27298
rect 26910 27246 26962 27298
rect 26962 27246 26964 27298
rect 26908 27244 26964 27246
rect 27244 31666 27300 31668
rect 27244 31614 27246 31666
rect 27246 31614 27298 31666
rect 27298 31614 27300 31666
rect 27244 31612 27300 31614
rect 28252 33964 28308 34020
rect 29596 43538 29652 43540
rect 29596 43486 29598 43538
rect 29598 43486 29650 43538
rect 29650 43486 29652 43538
rect 29596 43484 29652 43486
rect 30828 44546 30884 44548
rect 30828 44494 30830 44546
rect 30830 44494 30882 44546
rect 30882 44494 30884 44546
rect 30828 44492 30884 44494
rect 30604 44156 30660 44212
rect 29932 43372 29988 43428
rect 29372 42924 29428 42980
rect 29260 42700 29316 42756
rect 29036 42476 29092 42532
rect 29260 42530 29316 42532
rect 29260 42478 29262 42530
rect 29262 42478 29314 42530
rect 29314 42478 29316 42530
rect 29260 42476 29316 42478
rect 29148 40626 29204 40628
rect 29148 40574 29150 40626
rect 29150 40574 29202 40626
rect 29202 40574 29204 40626
rect 29148 40572 29204 40574
rect 29148 40012 29204 40068
rect 29148 38444 29204 38500
rect 28476 37266 28532 37268
rect 28476 37214 28478 37266
rect 28478 37214 28530 37266
rect 28530 37214 28532 37266
rect 28476 37212 28532 37214
rect 28588 35084 28644 35140
rect 28588 34412 28644 34468
rect 28476 33628 28532 33684
rect 28588 33458 28644 33460
rect 28588 33406 28590 33458
rect 28590 33406 28642 33458
rect 28642 33406 28644 33458
rect 28588 33404 28644 33406
rect 28252 33234 28308 33236
rect 28252 33182 28254 33234
rect 28254 33182 28306 33234
rect 28306 33182 28308 33234
rect 28252 33180 28308 33182
rect 28364 32396 28420 32452
rect 27580 31724 27636 31780
rect 27804 31948 27860 32004
rect 27580 31554 27636 31556
rect 27580 31502 27582 31554
rect 27582 31502 27634 31554
rect 27634 31502 27636 31554
rect 27580 31500 27636 31502
rect 27356 31106 27412 31108
rect 27356 31054 27358 31106
rect 27358 31054 27410 31106
rect 27410 31054 27412 31106
rect 27356 31052 27412 31054
rect 27692 30156 27748 30212
rect 27692 29596 27748 29652
rect 27244 28588 27300 28644
rect 27580 27804 27636 27860
rect 27356 27244 27412 27300
rect 27468 27132 27524 27188
rect 26796 26348 26852 26404
rect 26796 25228 26852 25284
rect 26796 24780 26852 24836
rect 26460 20130 26516 20132
rect 26460 20078 26462 20130
rect 26462 20078 26514 20130
rect 26514 20078 26516 20130
rect 26460 20076 26516 20078
rect 26460 19068 26516 19124
rect 25452 11788 25508 11844
rect 25676 14306 25732 14308
rect 25676 14254 25678 14306
rect 25678 14254 25730 14306
rect 25730 14254 25732 14306
rect 25676 14252 25732 14254
rect 25676 11340 25732 11396
rect 25004 10108 25060 10164
rect 23100 9996 23156 10052
rect 22764 9772 22820 9828
rect 23548 9826 23604 9828
rect 23548 9774 23550 9826
rect 23550 9774 23602 9826
rect 23602 9774 23604 9826
rect 23548 9772 23604 9774
rect 24332 9826 24388 9828
rect 24332 9774 24334 9826
rect 24334 9774 24386 9826
rect 24386 9774 24388 9826
rect 24332 9772 24388 9774
rect 24444 9714 24500 9716
rect 24444 9662 24446 9714
rect 24446 9662 24498 9714
rect 24498 9662 24500 9714
rect 24444 9660 24500 9662
rect 25900 9660 25956 9716
rect 21308 9042 21364 9044
rect 21308 8990 21310 9042
rect 21310 8990 21362 9042
rect 21362 8990 21364 9042
rect 21308 8988 21364 8990
rect 20188 6636 20244 6692
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 21084 7644 21140 7700
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 17836 3500 17892 3556
rect 19180 3554 19236 3556
rect 19180 3502 19182 3554
rect 19182 3502 19234 3554
rect 19234 3502 19236 3554
rect 19180 3500 19236 3502
rect 20860 3612 20916 3668
rect 20076 3554 20132 3556
rect 20076 3502 20078 3554
rect 20078 3502 20130 3554
rect 20130 3502 20132 3554
rect 20076 3500 20132 3502
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22204 9154 22260 9156
rect 22204 9102 22206 9154
rect 22206 9102 22258 9154
rect 22258 9102 22260 9154
rect 22204 9100 22260 9102
rect 21868 8988 21924 9044
rect 21868 7698 21924 7700
rect 21868 7646 21870 7698
rect 21870 7646 21922 7698
rect 21922 7646 21924 7698
rect 21868 7644 21924 7646
rect 22652 8316 22708 8372
rect 23660 8370 23716 8372
rect 23660 8318 23662 8370
rect 23662 8318 23714 8370
rect 23714 8318 23716 8370
rect 23660 8316 23716 8318
rect 22988 8258 23044 8260
rect 22988 8206 22990 8258
rect 22990 8206 23042 8258
rect 23042 8206 23044 8258
rect 22988 8204 23044 8206
rect 23660 6690 23716 6692
rect 23660 6638 23662 6690
rect 23662 6638 23714 6690
rect 23714 6638 23716 6690
rect 23660 6636 23716 6638
rect 24220 6690 24276 6692
rect 24220 6638 24222 6690
rect 24222 6638 24274 6690
rect 24274 6638 24276 6690
rect 24220 6636 24276 6638
rect 22652 5180 22708 5236
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 24108 5234 24164 5236
rect 24108 5182 24110 5234
rect 24110 5182 24162 5234
rect 24162 5182 24164 5234
rect 24108 5180 24164 5182
rect 26796 19964 26852 20020
rect 27244 25282 27300 25284
rect 27244 25230 27246 25282
rect 27246 25230 27298 25282
rect 27298 25230 27300 25282
rect 27244 25228 27300 25230
rect 27580 23884 27636 23940
rect 27692 23100 27748 23156
rect 27468 22092 27524 22148
rect 27020 20130 27076 20132
rect 27020 20078 27022 20130
rect 27022 20078 27074 20130
rect 27074 20078 27076 20130
rect 27020 20076 27076 20078
rect 28364 32172 28420 32228
rect 27916 28588 27972 28644
rect 28140 30994 28196 30996
rect 28140 30942 28142 30994
rect 28142 30942 28194 30994
rect 28194 30942 28196 30994
rect 28140 30940 28196 30942
rect 30492 41356 30548 41412
rect 30156 39730 30212 39732
rect 30156 39678 30158 39730
rect 30158 39678 30210 39730
rect 30210 39678 30212 39730
rect 30156 39676 30212 39678
rect 29484 39618 29540 39620
rect 29484 39566 29486 39618
rect 29486 39566 29538 39618
rect 29538 39566 29540 39618
rect 29484 39564 29540 39566
rect 29372 39004 29428 39060
rect 29372 37490 29428 37492
rect 29372 37438 29374 37490
rect 29374 37438 29426 37490
rect 29426 37438 29428 37490
rect 29372 37436 29428 37438
rect 29932 37266 29988 37268
rect 29932 37214 29934 37266
rect 29934 37214 29986 37266
rect 29986 37214 29988 37266
rect 29932 37212 29988 37214
rect 28700 32172 28756 32228
rect 30044 35084 30100 35140
rect 29820 34972 29876 35028
rect 29148 34802 29204 34804
rect 29148 34750 29150 34802
rect 29150 34750 29202 34802
rect 29202 34750 29204 34802
rect 29148 34748 29204 34750
rect 29708 34802 29764 34804
rect 29708 34750 29710 34802
rect 29710 34750 29762 34802
rect 29762 34750 29764 34802
rect 29708 34748 29764 34750
rect 29820 34412 29876 34468
rect 29148 33516 29204 33572
rect 29036 33180 29092 33236
rect 29484 33740 29540 33796
rect 29372 33346 29428 33348
rect 29372 33294 29374 33346
rect 29374 33294 29426 33346
rect 29426 33294 29428 33346
rect 29372 33292 29428 33294
rect 28588 30994 28644 30996
rect 28588 30942 28590 30994
rect 28590 30942 28642 30994
rect 28642 30942 28644 30994
rect 28588 30940 28644 30942
rect 28476 30268 28532 30324
rect 28476 29596 28532 29652
rect 28028 23100 28084 23156
rect 27132 19010 27188 19012
rect 27132 18958 27134 19010
rect 27134 18958 27186 19010
rect 27186 18958 27188 19010
rect 27132 18956 27188 18958
rect 26908 17836 26964 17892
rect 26796 15596 26852 15652
rect 26460 15202 26516 15204
rect 26460 15150 26462 15202
rect 26462 15150 26514 15202
rect 26514 15150 26516 15202
rect 26460 15148 26516 15150
rect 27132 14642 27188 14644
rect 27132 14590 27134 14642
rect 27134 14590 27186 14642
rect 27186 14590 27188 14642
rect 27132 14588 27188 14590
rect 26684 14306 26740 14308
rect 26684 14254 26686 14306
rect 26686 14254 26738 14306
rect 26738 14254 26740 14306
rect 26684 14252 26740 14254
rect 26348 13468 26404 13524
rect 26460 14140 26516 14196
rect 27244 14140 27300 14196
rect 27244 12850 27300 12852
rect 27244 12798 27246 12850
rect 27246 12798 27298 12850
rect 27298 12798 27300 12850
rect 27244 12796 27300 12798
rect 26348 11788 26404 11844
rect 26236 10834 26292 10836
rect 26236 10782 26238 10834
rect 26238 10782 26290 10834
rect 26290 10782 26292 10834
rect 26236 10780 26292 10782
rect 26236 8876 26292 8932
rect 26796 11788 26852 11844
rect 26908 11116 26964 11172
rect 27580 18956 27636 19012
rect 27468 17836 27524 17892
rect 27580 17554 27636 17556
rect 27580 17502 27582 17554
rect 27582 17502 27634 17554
rect 27634 17502 27636 17554
rect 27580 17500 27636 17502
rect 28252 23154 28308 23156
rect 28252 23102 28254 23154
rect 28254 23102 28306 23154
rect 28306 23102 28308 23154
rect 28252 23100 28308 23102
rect 28140 17500 28196 17556
rect 27804 15596 27860 15652
rect 27580 14140 27636 14196
rect 27916 15148 27972 15204
rect 28028 15260 28084 15316
rect 28588 24050 28644 24052
rect 28588 23998 28590 24050
rect 28590 23998 28642 24050
rect 28642 23998 28644 24050
rect 28588 23996 28644 23998
rect 29148 32060 29204 32116
rect 29036 31612 29092 31668
rect 29372 27692 29428 27748
rect 29484 26236 29540 26292
rect 29148 23996 29204 24052
rect 29484 23938 29540 23940
rect 29484 23886 29486 23938
rect 29486 23886 29538 23938
rect 29538 23886 29540 23938
rect 29484 23884 29540 23886
rect 30492 35196 30548 35252
rect 31612 43650 31668 43652
rect 31612 43598 31614 43650
rect 31614 43598 31666 43650
rect 31666 43598 31668 43650
rect 31612 43596 31668 43598
rect 31276 43538 31332 43540
rect 31276 43486 31278 43538
rect 31278 43486 31330 43538
rect 31330 43486 31332 43538
rect 31276 43484 31332 43486
rect 31164 41858 31220 41860
rect 31164 41806 31166 41858
rect 31166 41806 31218 41858
rect 31218 41806 31220 41858
rect 31164 41804 31220 41806
rect 30716 40908 30772 40964
rect 33180 46114 33236 46116
rect 33180 46062 33182 46114
rect 33182 46062 33234 46114
rect 33234 46062 33236 46114
rect 33180 46060 33236 46062
rect 33628 46060 33684 46116
rect 32284 44940 32340 44996
rect 33068 45836 33124 45892
rect 31724 40236 31780 40292
rect 32508 41804 32564 41860
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35980 45890 36036 45892
rect 35980 45838 35982 45890
rect 35982 45838 36034 45890
rect 36034 45838 36036 45890
rect 35980 45836 36036 45838
rect 34972 45276 35028 45332
rect 34412 45052 34468 45108
rect 33292 44994 33348 44996
rect 33292 44942 33294 44994
rect 33294 44942 33346 44994
rect 33346 44942 33348 44994
rect 33292 44940 33348 44942
rect 33404 44210 33460 44212
rect 33404 44158 33406 44210
rect 33406 44158 33458 44210
rect 33458 44158 33460 44210
rect 33404 44156 33460 44158
rect 33740 44210 33796 44212
rect 33740 44158 33742 44210
rect 33742 44158 33794 44210
rect 33794 44158 33796 44210
rect 33740 44156 33796 44158
rect 33404 43708 33460 43764
rect 33180 43538 33236 43540
rect 33180 43486 33182 43538
rect 33182 43486 33234 43538
rect 33234 43486 33236 43538
rect 33180 43484 33236 43486
rect 32732 41356 32788 41412
rect 30716 40124 30772 40180
rect 31500 40124 31556 40180
rect 30828 39900 30884 39956
rect 30828 39004 30884 39060
rect 30716 38722 30772 38724
rect 30716 38670 30718 38722
rect 30718 38670 30770 38722
rect 30770 38670 30772 38722
rect 30716 38668 30772 38670
rect 32284 39788 32340 39844
rect 32732 39618 32788 39620
rect 32732 39566 32734 39618
rect 32734 39566 32786 39618
rect 32786 39566 32788 39618
rect 32732 39564 32788 39566
rect 32508 39058 32564 39060
rect 32508 39006 32510 39058
rect 32510 39006 32562 39058
rect 32562 39006 32564 39058
rect 32508 39004 32564 39006
rect 32508 37490 32564 37492
rect 32508 37438 32510 37490
rect 32510 37438 32562 37490
rect 32562 37438 32564 37490
rect 32508 37436 32564 37438
rect 33404 39116 33460 39172
rect 35196 45106 35252 45108
rect 35196 45054 35198 45106
rect 35198 45054 35250 45106
rect 35250 45054 35252 45106
rect 35196 45052 35252 45054
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35644 44268 35700 44324
rect 36988 46114 37044 46116
rect 36988 46062 36990 46114
rect 36990 46062 37042 46114
rect 37042 46062 37044 46114
rect 36988 46060 37044 46062
rect 37660 46060 37716 46116
rect 36988 45330 37044 45332
rect 36988 45278 36990 45330
rect 36990 45278 37042 45330
rect 37042 45278 37044 45330
rect 36988 45276 37044 45278
rect 36316 44492 36372 44548
rect 37996 44546 38052 44548
rect 37996 44494 37998 44546
rect 37998 44494 38050 44546
rect 38050 44494 38052 44546
rect 37996 44492 38052 44494
rect 39788 45500 39844 45556
rect 40796 46114 40852 46116
rect 40796 46062 40798 46114
rect 40798 46062 40850 46114
rect 40850 46062 40852 46114
rect 40796 46060 40852 46062
rect 41692 46060 41748 46116
rect 40348 45276 40404 45332
rect 41916 45330 41972 45332
rect 41916 45278 41918 45330
rect 41918 45278 41970 45330
rect 41970 45278 41972 45330
rect 41916 45276 41972 45278
rect 43036 45276 43092 45332
rect 39004 44492 39060 44548
rect 40908 44546 40964 44548
rect 40908 44494 40910 44546
rect 40910 44494 40962 44546
rect 40962 44494 40964 44546
rect 40908 44492 40964 44494
rect 36988 44322 37044 44324
rect 36988 44270 36990 44322
rect 36990 44270 37042 44322
rect 37042 44270 37044 44322
rect 36988 44268 37044 44270
rect 39900 44156 39956 44212
rect 35980 43708 36036 43764
rect 37324 43484 37380 43540
rect 34188 40236 34244 40292
rect 33292 38722 33348 38724
rect 33292 38670 33294 38722
rect 33294 38670 33346 38722
rect 33346 38670 33348 38722
rect 33292 38668 33348 38670
rect 33180 37436 33236 37492
rect 32172 36204 32228 36260
rect 32508 35586 32564 35588
rect 32508 35534 32510 35586
rect 32510 35534 32562 35586
rect 32562 35534 32564 35586
rect 32508 35532 32564 35534
rect 30268 35026 30324 35028
rect 30268 34974 30270 35026
rect 30270 34974 30322 35026
rect 30322 34974 30324 35026
rect 30268 34972 30324 34974
rect 29708 33234 29764 33236
rect 29708 33182 29710 33234
rect 29710 33182 29762 33234
rect 29762 33182 29764 33234
rect 29708 33180 29764 33182
rect 30268 34748 30324 34804
rect 29708 32060 29764 32116
rect 29708 28588 29764 28644
rect 29932 27746 29988 27748
rect 29932 27694 29934 27746
rect 29934 27694 29986 27746
rect 29986 27694 29988 27746
rect 29932 27692 29988 27694
rect 30380 33234 30436 33236
rect 30380 33182 30382 33234
rect 30382 33182 30434 33234
rect 30434 33182 30436 33234
rect 30380 33180 30436 33182
rect 30828 35084 30884 35140
rect 30380 31052 30436 31108
rect 30716 30098 30772 30100
rect 30716 30046 30718 30098
rect 30718 30046 30770 30098
rect 30770 30046 30772 30098
rect 30716 30044 30772 30046
rect 30268 27804 30324 27860
rect 30156 27468 30212 27524
rect 31164 30210 31220 30212
rect 31164 30158 31166 30210
rect 31166 30158 31218 30210
rect 31218 30158 31220 30210
rect 31164 30156 31220 30158
rect 31836 30268 31892 30324
rect 30940 29650 30996 29652
rect 30940 29598 30942 29650
rect 30942 29598 30994 29650
rect 30994 29598 30996 29650
rect 30940 29596 30996 29598
rect 31276 29484 31332 29540
rect 32732 35026 32788 35028
rect 32732 34974 32734 35026
rect 32734 34974 32786 35026
rect 32786 34974 32788 35026
rect 32732 34972 32788 34974
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34972 39788 35028 39844
rect 34524 38946 34580 38948
rect 34524 38894 34526 38946
rect 34526 38894 34578 38946
rect 34578 38894 34580 38946
rect 34524 38892 34580 38894
rect 34300 38722 34356 38724
rect 34300 38670 34302 38722
rect 34302 38670 34354 38722
rect 34354 38670 34356 38722
rect 34300 38668 34356 38670
rect 35532 39788 35588 39844
rect 33740 37378 33796 37380
rect 33740 37326 33742 37378
rect 33742 37326 33794 37378
rect 33794 37326 33796 37378
rect 33740 37324 33796 37326
rect 33964 37154 34020 37156
rect 33964 37102 33966 37154
rect 33966 37102 34018 37154
rect 34018 37102 34020 37154
rect 33964 37100 34020 37102
rect 33740 36988 33796 37044
rect 33852 35586 33908 35588
rect 33852 35534 33854 35586
rect 33854 35534 33906 35586
rect 33906 35534 33908 35586
rect 33852 35532 33908 35534
rect 33516 33964 33572 34020
rect 31948 28364 32004 28420
rect 32172 28476 32228 28532
rect 31836 27692 31892 27748
rect 30492 24722 30548 24724
rect 30492 24670 30494 24722
rect 30494 24670 30546 24722
rect 30546 24670 30548 24722
rect 30492 24668 30548 24670
rect 30828 23996 30884 24052
rect 29596 23772 29652 23828
rect 28812 22988 28868 23044
rect 29708 23042 29764 23044
rect 29708 22990 29710 23042
rect 29710 22990 29762 23042
rect 29762 22990 29764 23042
rect 29708 22988 29764 22990
rect 30268 22988 30324 23044
rect 31948 27186 32004 27188
rect 31948 27134 31950 27186
rect 31950 27134 32002 27186
rect 32002 27134 32004 27186
rect 31948 27132 32004 27134
rect 31612 26236 31668 26292
rect 31052 24722 31108 24724
rect 31052 24670 31054 24722
rect 31054 24670 31106 24722
rect 31106 24670 31108 24722
rect 31052 24668 31108 24670
rect 31500 23938 31556 23940
rect 31500 23886 31502 23938
rect 31502 23886 31554 23938
rect 31554 23886 31556 23938
rect 31500 23884 31556 23886
rect 29596 22092 29652 22148
rect 29372 20802 29428 20804
rect 29372 20750 29374 20802
rect 29374 20750 29426 20802
rect 29426 20750 29428 20802
rect 29372 20748 29428 20750
rect 30044 22092 30100 22148
rect 30044 21868 30100 21924
rect 29932 20802 29988 20804
rect 29932 20750 29934 20802
rect 29934 20750 29986 20802
rect 29986 20750 29988 20802
rect 29932 20748 29988 20750
rect 29708 19180 29764 19236
rect 28588 17442 28644 17444
rect 28588 17390 28590 17442
rect 28590 17390 28642 17442
rect 28642 17390 28644 17442
rect 28588 17388 28644 17390
rect 28588 15314 28644 15316
rect 28588 15262 28590 15314
rect 28590 15262 28642 15314
rect 28642 15262 28644 15314
rect 28588 15260 28644 15262
rect 27916 13804 27972 13860
rect 27356 12124 27412 12180
rect 27804 13356 27860 13412
rect 27692 12796 27748 12852
rect 27916 12178 27972 12180
rect 27916 12126 27918 12178
rect 27918 12126 27970 12178
rect 27970 12126 27972 12178
rect 27916 12124 27972 12126
rect 27244 10780 27300 10836
rect 26908 9996 26964 10052
rect 27132 8930 27188 8932
rect 27132 8878 27134 8930
rect 27134 8878 27186 8930
rect 27186 8878 27188 8930
rect 27132 8876 27188 8878
rect 28588 14252 28644 14308
rect 28476 13858 28532 13860
rect 28476 13806 28478 13858
rect 28478 13806 28530 13858
rect 28530 13806 28532 13858
rect 28476 13804 28532 13806
rect 28588 13074 28644 13076
rect 28588 13022 28590 13074
rect 28590 13022 28642 13074
rect 28642 13022 28644 13074
rect 28588 13020 28644 13022
rect 28588 12178 28644 12180
rect 28588 12126 28590 12178
rect 28590 12126 28642 12178
rect 28642 12126 28644 12178
rect 28588 12124 28644 12126
rect 26348 8258 26404 8260
rect 26348 8206 26350 8258
rect 26350 8206 26402 8258
rect 26402 8206 26404 8258
rect 26348 8204 26404 8206
rect 29036 18060 29092 18116
rect 29372 17500 29428 17556
rect 29148 17106 29204 17108
rect 29148 17054 29150 17106
rect 29150 17054 29202 17106
rect 29202 17054 29204 17106
rect 29148 17052 29204 17054
rect 30828 23100 30884 23156
rect 30156 20690 30212 20692
rect 30156 20638 30158 20690
rect 30158 20638 30210 20690
rect 30210 20638 30212 20690
rect 30156 20636 30212 20638
rect 31724 21756 31780 21812
rect 32060 21532 32116 21588
rect 30268 20076 30324 20132
rect 30268 19740 30324 19796
rect 30828 20188 30884 20244
rect 31836 20188 31892 20244
rect 30716 20130 30772 20132
rect 30716 20078 30718 20130
rect 30718 20078 30770 20130
rect 30770 20078 30772 20130
rect 30716 20076 30772 20078
rect 30828 19740 30884 19796
rect 30604 19234 30660 19236
rect 30604 19182 30606 19234
rect 30606 19182 30658 19234
rect 30658 19182 30660 19234
rect 30604 19180 30660 19182
rect 30492 18450 30548 18452
rect 30492 18398 30494 18450
rect 30494 18398 30546 18450
rect 30546 18398 30548 18450
rect 30492 18396 30548 18398
rect 29820 18060 29876 18116
rect 30716 19010 30772 19012
rect 30716 18958 30718 19010
rect 30718 18958 30770 19010
rect 30770 18958 30772 19010
rect 30716 18956 30772 18958
rect 30380 17500 30436 17556
rect 30716 17554 30772 17556
rect 30716 17502 30718 17554
rect 30718 17502 30770 17554
rect 30770 17502 30772 17554
rect 30716 17500 30772 17502
rect 30604 17388 30660 17444
rect 30156 16268 30212 16324
rect 29596 16156 29652 16212
rect 29932 15708 29988 15764
rect 30268 15538 30324 15540
rect 30268 15486 30270 15538
rect 30270 15486 30322 15538
rect 30322 15486 30324 15538
rect 30268 15484 30324 15486
rect 29260 15148 29316 15204
rect 28924 14476 28980 14532
rect 28924 13970 28980 13972
rect 28924 13918 28926 13970
rect 28926 13918 28978 13970
rect 28978 13918 28980 13970
rect 28924 13916 28980 13918
rect 30156 15148 30212 15204
rect 30156 14530 30212 14532
rect 30156 14478 30158 14530
rect 30158 14478 30210 14530
rect 30210 14478 30212 14530
rect 30156 14476 30212 14478
rect 29708 13468 29764 13524
rect 29372 13020 29428 13076
rect 30044 12962 30100 12964
rect 30044 12910 30046 12962
rect 30046 12910 30098 12962
rect 30098 12910 30100 12962
rect 30044 12908 30100 12910
rect 29260 12178 29316 12180
rect 29260 12126 29262 12178
rect 29262 12126 29314 12178
rect 29314 12126 29316 12178
rect 29260 12124 29316 12126
rect 30044 12572 30100 12628
rect 29148 11676 29204 11732
rect 29148 10444 29204 10500
rect 29708 10498 29764 10500
rect 29708 10446 29710 10498
rect 29710 10446 29762 10498
rect 29762 10446 29764 10498
rect 29708 10444 29764 10446
rect 31724 19740 31780 19796
rect 31388 18956 31444 19012
rect 31948 19852 32004 19908
rect 32172 19292 32228 19348
rect 31388 18338 31444 18340
rect 31388 18286 31390 18338
rect 31390 18286 31442 18338
rect 31442 18286 31444 18338
rect 31388 18284 31444 18286
rect 31836 18338 31892 18340
rect 31836 18286 31838 18338
rect 31838 18286 31890 18338
rect 31890 18286 31892 18338
rect 31836 18284 31892 18286
rect 30940 17164 30996 17220
rect 30940 15932 30996 15988
rect 30716 15820 30772 15876
rect 31500 17164 31556 17220
rect 31612 16604 31668 16660
rect 31724 16940 31780 16996
rect 31164 16044 31220 16100
rect 31500 16044 31556 16100
rect 31388 15986 31444 15988
rect 31388 15934 31390 15986
rect 31390 15934 31442 15986
rect 31442 15934 31444 15986
rect 31388 15932 31444 15934
rect 32060 16156 32116 16212
rect 31164 15874 31220 15876
rect 31164 15822 31166 15874
rect 31166 15822 31218 15874
rect 31218 15822 31220 15874
rect 31164 15820 31220 15822
rect 30716 14252 30772 14308
rect 30828 13858 30884 13860
rect 30828 13806 30830 13858
rect 30830 13806 30882 13858
rect 30882 13806 30884 13858
rect 30828 13804 30884 13806
rect 30604 13244 30660 13300
rect 30268 12908 30324 12964
rect 30492 12738 30548 12740
rect 30492 12686 30494 12738
rect 30494 12686 30546 12738
rect 30546 12686 30548 12738
rect 30492 12684 30548 12686
rect 30380 12178 30436 12180
rect 30380 12126 30382 12178
rect 30382 12126 30434 12178
rect 30434 12126 30436 12178
rect 30380 12124 30436 12126
rect 30156 11900 30212 11956
rect 31724 15538 31780 15540
rect 31724 15486 31726 15538
rect 31726 15486 31778 15538
rect 31778 15486 31780 15538
rect 31724 15484 31780 15486
rect 31612 13804 31668 13860
rect 31052 13244 31108 13300
rect 31276 13020 31332 13076
rect 31388 13468 31444 13524
rect 31052 12572 31108 12628
rect 30604 11452 30660 11508
rect 30940 11676 30996 11732
rect 30268 9548 30324 9604
rect 31500 12738 31556 12740
rect 31500 12686 31502 12738
rect 31502 12686 31554 12738
rect 31554 12686 31556 12738
rect 31500 12684 31556 12686
rect 31948 11788 32004 11844
rect 31612 11452 31668 11508
rect 32172 9602 32228 9604
rect 32172 9550 32174 9602
rect 32174 9550 32226 9602
rect 32226 9550 32228 9602
rect 32172 9548 32228 9550
rect 33628 31948 33684 32004
rect 32732 31164 32788 31220
rect 32396 28364 32452 28420
rect 32508 27746 32564 27748
rect 32508 27694 32510 27746
rect 32510 27694 32562 27746
rect 32562 27694 32564 27746
rect 32508 27692 32564 27694
rect 32396 27132 32452 27188
rect 33068 30156 33124 30212
rect 33628 31612 33684 31668
rect 33180 29148 33236 29204
rect 33852 32060 33908 32116
rect 34076 33180 34132 33236
rect 33740 31218 33796 31220
rect 33740 31166 33742 31218
rect 33742 31166 33794 31218
rect 33794 31166 33796 31218
rect 33740 31164 33796 31166
rect 33852 31724 33908 31780
rect 33852 31052 33908 31108
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34860 37378 34916 37380
rect 34860 37326 34862 37378
rect 34862 37326 34914 37378
rect 34914 37326 34916 37378
rect 34860 37324 34916 37326
rect 35420 37154 35476 37156
rect 35420 37102 35422 37154
rect 35422 37102 35474 37154
rect 35474 37102 35476 37154
rect 35420 37100 35476 37102
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34748 36204 34804 36260
rect 34524 35084 34580 35140
rect 35084 35532 35140 35588
rect 35532 35420 35588 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34524 32956 34580 33012
rect 34412 32732 34468 32788
rect 34524 32620 34580 32676
rect 34188 31612 34244 31668
rect 34076 31500 34132 31556
rect 34188 31218 34244 31220
rect 34188 31166 34190 31218
rect 34190 31166 34242 31218
rect 34242 31166 34244 31218
rect 34188 31164 34244 31166
rect 34076 30940 34132 30996
rect 34188 30492 34244 30548
rect 33628 28028 33684 28084
rect 33852 27746 33908 27748
rect 33852 27694 33854 27746
rect 33854 27694 33906 27746
rect 33906 27694 33908 27746
rect 33852 27692 33908 27694
rect 34412 30156 34468 30212
rect 35532 33852 35588 33908
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35980 39618 36036 39620
rect 35980 39566 35982 39618
rect 35982 39566 36034 39618
rect 36034 39566 36036 39618
rect 35980 39564 36036 39566
rect 36092 38946 36148 38948
rect 36092 38894 36094 38946
rect 36094 38894 36146 38946
rect 36146 38894 36148 38946
rect 36092 38892 36148 38894
rect 36652 38722 36708 38724
rect 36652 38670 36654 38722
rect 36654 38670 36706 38722
rect 36706 38670 36708 38722
rect 36652 38668 36708 38670
rect 35868 37100 35924 37156
rect 35980 35586 36036 35588
rect 35980 35534 35982 35586
rect 35982 35534 36034 35586
rect 36034 35534 36036 35586
rect 35980 35532 36036 35534
rect 35532 33458 35588 33460
rect 35532 33406 35534 33458
rect 35534 33406 35586 33458
rect 35586 33406 35588 33458
rect 35532 33404 35588 33406
rect 34860 32956 34916 33012
rect 35868 33346 35924 33348
rect 35868 33294 35870 33346
rect 35870 33294 35922 33346
rect 35922 33294 35924 33346
rect 35868 33292 35924 33294
rect 35756 33234 35812 33236
rect 35756 33182 35758 33234
rect 35758 33182 35810 33234
rect 35810 33182 35812 33234
rect 35756 33180 35812 33182
rect 34860 32674 34916 32676
rect 34860 32622 34862 32674
rect 34862 32622 34914 32674
rect 34914 32622 34916 32674
rect 34860 32620 34916 32622
rect 35420 32284 35476 32340
rect 35756 32508 35812 32564
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 34748 31948 34804 32004
rect 34860 31106 34916 31108
rect 34860 31054 34862 31106
rect 34862 31054 34914 31106
rect 34914 31054 34916 31106
rect 34860 31052 34916 31054
rect 37212 35420 37268 35476
rect 36092 35026 36148 35028
rect 36092 34974 36094 35026
rect 36094 34974 36146 35026
rect 36146 34974 36148 35026
rect 36092 34972 36148 34974
rect 36876 32732 36932 32788
rect 36428 32562 36484 32564
rect 36428 32510 36430 32562
rect 36430 32510 36482 32562
rect 36482 32510 36484 32562
rect 36428 32508 36484 32510
rect 36316 32450 36372 32452
rect 36316 32398 36318 32450
rect 36318 32398 36370 32450
rect 36370 32398 36372 32450
rect 36316 32396 36372 32398
rect 36876 32284 36932 32340
rect 36876 31948 36932 32004
rect 34748 30380 34804 30436
rect 34860 30828 34916 30884
rect 34636 29484 34692 29540
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35532 30268 35588 30324
rect 34412 27916 34468 27972
rect 32844 25788 32900 25844
rect 32396 25564 32452 25620
rect 33516 26796 33572 26852
rect 35756 30098 35812 30100
rect 35756 30046 35758 30098
rect 35758 30046 35810 30098
rect 35810 30046 35812 30098
rect 35756 30044 35812 30046
rect 35420 29484 35476 29540
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34860 28588 34916 28644
rect 34748 28530 34804 28532
rect 34748 28478 34750 28530
rect 34750 28478 34802 28530
rect 34802 28478 34804 28530
rect 34748 28476 34804 28478
rect 34972 27692 35028 27748
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 33292 25564 33348 25620
rect 33404 26124 33460 26180
rect 33516 25900 33572 25956
rect 33628 25788 33684 25844
rect 33404 25340 33460 25396
rect 34524 26684 34580 26740
rect 34412 26460 34468 26516
rect 34300 25788 34356 25844
rect 34188 25394 34244 25396
rect 34188 25342 34190 25394
rect 34190 25342 34242 25394
rect 34242 25342 34244 25394
rect 34188 25340 34244 25342
rect 33852 24780 33908 24836
rect 34300 25004 34356 25060
rect 33180 22988 33236 23044
rect 33628 24444 33684 24500
rect 33068 20690 33124 20692
rect 33068 20638 33070 20690
rect 33070 20638 33122 20690
rect 33122 20638 33124 20690
rect 33068 20636 33124 20638
rect 32844 19292 32900 19348
rect 32396 15596 32452 15652
rect 32284 9100 32340 9156
rect 32732 18284 32788 18340
rect 33852 20860 33908 20916
rect 33628 18956 33684 19012
rect 33292 18284 33348 18340
rect 33180 17164 33236 17220
rect 32732 16604 32788 16660
rect 33068 15932 33124 15988
rect 33180 15484 33236 15540
rect 33740 17164 33796 17220
rect 33404 16882 33460 16884
rect 33404 16830 33406 16882
rect 33406 16830 33458 16882
rect 33458 16830 33460 16882
rect 33404 16828 33460 16830
rect 33292 14476 33348 14532
rect 33628 16268 33684 16324
rect 32732 13074 32788 13076
rect 32732 13022 32734 13074
rect 32734 13022 32786 13074
rect 32786 13022 32788 13074
rect 32732 13020 32788 13022
rect 32732 11116 32788 11172
rect 32732 10444 32788 10500
rect 31164 7644 31220 7700
rect 28700 6636 28756 6692
rect 28252 5964 28308 6020
rect 29036 5964 29092 6020
rect 26908 4060 26964 4116
rect 26124 3500 26180 3556
rect 28140 4114 28196 4116
rect 28140 4062 28142 4114
rect 28142 4062 28194 4114
rect 28194 4062 28196 4114
rect 28140 4060 28196 4062
rect 27244 3554 27300 3556
rect 27244 3502 27246 3554
rect 27246 3502 27298 3554
rect 27298 3502 27300 3554
rect 27244 3500 27300 3502
rect 28476 3554 28532 3556
rect 28476 3502 28478 3554
rect 28478 3502 28530 3554
rect 28530 3502 28532 3554
rect 28476 3500 28532 3502
rect 32956 4060 33012 4116
rect 32620 3554 32676 3556
rect 32620 3502 32622 3554
rect 32622 3502 32674 3554
rect 32674 3502 32676 3554
rect 32620 3500 32676 3502
rect 28924 3388 28980 3444
rect 30044 3388 30100 3444
rect 30940 3388 30996 3444
rect 34636 25900 34692 25956
rect 34412 24892 34468 24948
rect 34524 25340 34580 25396
rect 35980 30716 36036 30772
rect 36988 31836 37044 31892
rect 39788 42642 39844 42644
rect 39788 42590 39790 42642
rect 39790 42590 39842 42642
rect 39842 42590 39844 42642
rect 39788 42588 39844 42590
rect 40796 42642 40852 42644
rect 40796 42590 40798 42642
rect 40798 42590 40850 42642
rect 40850 42590 40852 42642
rect 40796 42588 40852 42590
rect 39228 42476 39284 42532
rect 39116 37938 39172 37940
rect 39116 37886 39118 37938
rect 39118 37886 39170 37938
rect 39170 37886 39172 37938
rect 39116 37884 39172 37886
rect 39004 37772 39060 37828
rect 38668 35756 38724 35812
rect 36988 31218 37044 31220
rect 36988 31166 36990 31218
rect 36990 31166 37042 31218
rect 37042 31166 37044 31218
rect 36988 31164 37044 31166
rect 37100 31554 37156 31556
rect 37100 31502 37102 31554
rect 37102 31502 37154 31554
rect 37154 31502 37156 31554
rect 37100 31500 37156 31502
rect 36540 30994 36596 30996
rect 36540 30942 36542 30994
rect 36542 30942 36594 30994
rect 36594 30942 36596 30994
rect 36540 30940 36596 30942
rect 36988 30770 37044 30772
rect 36988 30718 36990 30770
rect 36990 30718 37042 30770
rect 37042 30718 37044 30770
rect 36988 30716 37044 30718
rect 35980 29260 36036 29316
rect 35980 27746 36036 27748
rect 35980 27694 35982 27746
rect 35982 27694 36034 27746
rect 36034 27694 36036 27746
rect 35980 27692 36036 27694
rect 35532 27074 35588 27076
rect 35532 27022 35534 27074
rect 35534 27022 35586 27074
rect 35586 27022 35588 27074
rect 35532 27020 35588 27022
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35084 25564 35140 25620
rect 34972 25452 35028 25508
rect 34860 25394 34916 25396
rect 34860 25342 34862 25394
rect 34862 25342 34914 25394
rect 34914 25342 34916 25394
rect 34860 25340 34916 25342
rect 34748 24780 34804 24836
rect 34076 24610 34132 24612
rect 34076 24558 34078 24610
rect 34078 24558 34130 24610
rect 34130 24558 34132 24610
rect 34076 24556 34132 24558
rect 34412 24220 34468 24276
rect 34076 24108 34132 24164
rect 34188 22092 34244 22148
rect 34412 21810 34468 21812
rect 34412 21758 34414 21810
rect 34414 21758 34466 21810
rect 34466 21758 34468 21810
rect 34412 21756 34468 21758
rect 34860 24556 34916 24612
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21810 35252 21812
rect 35196 21758 35198 21810
rect 35198 21758 35250 21810
rect 35250 21758 35252 21810
rect 35196 21756 35252 21758
rect 34748 21532 34804 21588
rect 35420 21532 35476 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34972 20914 35028 20916
rect 34972 20862 34974 20914
rect 34974 20862 35026 20914
rect 35026 20862 35028 20914
rect 34972 20860 35028 20862
rect 35084 20076 35140 20132
rect 34860 19852 34916 19908
rect 35532 20130 35588 20132
rect 35532 20078 35534 20130
rect 35534 20078 35586 20130
rect 35586 20078 35588 20130
rect 35532 20076 35588 20078
rect 35196 20018 35252 20020
rect 35196 19966 35198 20018
rect 35198 19966 35250 20018
rect 35250 19966 35252 20018
rect 35196 19964 35252 19966
rect 35420 19852 35476 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34636 19180 34692 19236
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34412 17500 34468 17556
rect 35420 17052 35476 17108
rect 35532 16994 35588 16996
rect 35532 16942 35534 16994
rect 35534 16942 35586 16994
rect 35586 16942 35588 16994
rect 35532 16940 35588 16942
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35532 16210 35588 16212
rect 35532 16158 35534 16210
rect 35534 16158 35586 16210
rect 35586 16158 35588 16210
rect 35532 16156 35588 16158
rect 34860 15820 34916 15876
rect 36316 27074 36372 27076
rect 36316 27022 36318 27074
rect 36318 27022 36370 27074
rect 36370 27022 36372 27074
rect 36316 27020 36372 27022
rect 35868 26684 35924 26740
rect 36204 26796 36260 26852
rect 38220 32450 38276 32452
rect 38220 32398 38222 32450
rect 38222 32398 38274 32450
rect 38274 32398 38276 32450
rect 38220 32396 38276 32398
rect 37436 31500 37492 31556
rect 37996 31218 38052 31220
rect 37996 31166 37998 31218
rect 37998 31166 38050 31218
rect 38050 31166 38052 31218
rect 37996 31164 38052 31166
rect 37548 30380 37604 30436
rect 37212 30156 37268 30212
rect 37100 29932 37156 29988
rect 38556 29986 38612 29988
rect 38556 29934 38558 29986
rect 38558 29934 38610 29986
rect 38610 29934 38612 29986
rect 38556 29932 38612 29934
rect 36428 26460 36484 26516
rect 35756 25618 35812 25620
rect 35756 25566 35758 25618
rect 35758 25566 35810 25618
rect 35810 25566 35812 25618
rect 35756 25564 35812 25566
rect 36316 25340 36372 25396
rect 36428 24668 36484 24724
rect 39004 35756 39060 35812
rect 38892 33458 38948 33460
rect 38892 33406 38894 33458
rect 38894 33406 38946 33458
rect 38946 33406 38948 33458
rect 38892 33404 38948 33406
rect 38892 29932 38948 29988
rect 38780 28700 38836 28756
rect 37100 26796 37156 26852
rect 38556 26796 38612 26852
rect 36876 26178 36932 26180
rect 36876 26126 36878 26178
rect 36878 26126 36930 26178
rect 36930 26126 36932 26178
rect 36876 26124 36932 26126
rect 37996 26178 38052 26180
rect 37996 26126 37998 26178
rect 37998 26126 38050 26178
rect 38050 26126 38052 26178
rect 37996 26124 38052 26126
rect 36876 24668 36932 24724
rect 36652 24498 36708 24500
rect 36652 24446 36654 24498
rect 36654 24446 36706 24498
rect 36706 24446 36708 24498
rect 36652 24444 36708 24446
rect 37772 24444 37828 24500
rect 36428 23884 36484 23940
rect 37100 23938 37156 23940
rect 37100 23886 37102 23938
rect 37102 23886 37154 23938
rect 37154 23886 37156 23938
rect 37100 23884 37156 23886
rect 37884 23884 37940 23940
rect 35756 20578 35812 20580
rect 35756 20526 35758 20578
rect 35758 20526 35810 20578
rect 35810 20526 35812 20578
rect 35756 20524 35812 20526
rect 36652 20524 36708 20580
rect 35756 20188 35812 20244
rect 36540 20018 36596 20020
rect 36540 19966 36542 20018
rect 36542 19966 36594 20018
rect 36594 19966 36596 20018
rect 36540 19964 36596 19966
rect 36428 19906 36484 19908
rect 36428 19854 36430 19906
rect 36430 19854 36482 19906
rect 36482 19854 36484 19906
rect 36428 19852 36484 19854
rect 35980 19180 36036 19236
rect 35868 19010 35924 19012
rect 35868 18958 35870 19010
rect 35870 18958 35922 19010
rect 35922 18958 35924 19010
rect 35868 18956 35924 18958
rect 35868 18396 35924 18452
rect 36428 19234 36484 19236
rect 36428 19182 36430 19234
rect 36430 19182 36482 19234
rect 36482 19182 36484 19234
rect 36428 19180 36484 19182
rect 36316 19010 36372 19012
rect 36316 18958 36318 19010
rect 36318 18958 36370 19010
rect 36370 18958 36372 19010
rect 36316 18956 36372 18958
rect 35868 17388 35924 17444
rect 35756 15372 35812 15428
rect 36092 17442 36148 17444
rect 36092 17390 36094 17442
rect 36094 17390 36146 17442
rect 36146 17390 36148 17442
rect 36092 17388 36148 17390
rect 37212 20860 37268 20916
rect 37212 20188 37268 20244
rect 37884 20860 37940 20916
rect 37436 20690 37492 20692
rect 37436 20638 37438 20690
rect 37438 20638 37490 20690
rect 37490 20638 37492 20690
rect 37436 20636 37492 20638
rect 37884 20300 37940 20356
rect 37212 19292 37268 19348
rect 36988 19234 37044 19236
rect 36988 19182 36990 19234
rect 36990 19182 37042 19234
rect 37042 19182 37044 19234
rect 36988 19180 37044 19182
rect 37100 17442 37156 17444
rect 37100 17390 37102 17442
rect 37102 17390 37154 17442
rect 37154 17390 37156 17442
rect 37100 17388 37156 17390
rect 36428 17052 36484 17108
rect 36428 16882 36484 16884
rect 36428 16830 36430 16882
rect 36430 16830 36482 16882
rect 36482 16830 36484 16882
rect 36428 16828 36484 16830
rect 36316 16770 36372 16772
rect 36316 16718 36318 16770
rect 36318 16718 36370 16770
rect 36370 16718 36372 16770
rect 36316 16716 36372 16718
rect 37100 16268 37156 16324
rect 36316 16156 36372 16212
rect 35868 15260 35924 15316
rect 35980 15874 36036 15876
rect 35980 15822 35982 15874
rect 35982 15822 36034 15874
rect 36034 15822 36036 15874
rect 35980 15820 36036 15822
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35868 14252 35924 14308
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 34188 13020 34244 13076
rect 34860 13074 34916 13076
rect 34860 13022 34862 13074
rect 34862 13022 34914 13074
rect 34914 13022 34916 13074
rect 34860 13020 34916 13022
rect 33964 11676 34020 11732
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34524 11170 34580 11172
rect 34524 11118 34526 11170
rect 34526 11118 34578 11170
rect 34578 11118 34580 11170
rect 34524 11116 34580 11118
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 36988 16156 37044 16212
rect 37660 16156 37716 16212
rect 37772 16716 37828 16772
rect 37212 15820 37268 15876
rect 37100 15426 37156 15428
rect 37100 15374 37102 15426
rect 37102 15374 37154 15426
rect 37154 15374 37156 15426
rect 37100 15372 37156 15374
rect 35980 8876 36036 8932
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35980 4956 36036 5012
rect 34188 4114 34244 4116
rect 34188 4062 34190 4114
rect 34190 4062 34242 4114
rect 34242 4062 34244 4114
rect 34188 4060 34244 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 33628 3500 33684 3556
rect 33740 3442 33796 3444
rect 33740 3390 33742 3442
rect 33742 3390 33794 3442
rect 33794 3390 33796 3442
rect 33740 3388 33796 3390
rect 35532 3442 35588 3444
rect 35532 3390 35534 3442
rect 35534 3390 35586 3442
rect 35586 3390 35588 3442
rect 35532 3388 35588 3390
rect 36204 3388 36260 3444
rect 37996 19906 38052 19908
rect 37996 19854 37998 19906
rect 37998 19854 38050 19906
rect 38050 19854 38052 19906
rect 37996 19852 38052 19854
rect 38108 19346 38164 19348
rect 38108 19294 38110 19346
rect 38110 19294 38162 19346
rect 38162 19294 38164 19346
rect 38108 19292 38164 19294
rect 38892 25506 38948 25508
rect 38892 25454 38894 25506
rect 38894 25454 38946 25506
rect 38946 25454 38948 25506
rect 38892 25452 38948 25454
rect 39004 20690 39060 20692
rect 39004 20638 39006 20690
rect 39006 20638 39058 20690
rect 39058 20638 39060 20690
rect 39004 20636 39060 20638
rect 39116 20188 39172 20244
rect 40236 42530 40292 42532
rect 40236 42478 40238 42530
rect 40238 42478 40290 42530
rect 40290 42478 40292 42530
rect 40236 42476 40292 42478
rect 39788 41468 39844 41524
rect 39788 38050 39844 38052
rect 39788 37998 39790 38050
rect 39790 37998 39842 38050
rect 39842 37998 39844 38050
rect 39788 37996 39844 37998
rect 39340 37884 39396 37940
rect 39340 35084 39396 35140
rect 40908 42476 40964 42532
rect 41580 44380 41636 44436
rect 41916 44156 41972 44212
rect 42812 44210 42868 44212
rect 42812 44158 42814 44210
rect 42814 44158 42866 44210
rect 42866 44158 42868 44210
rect 42812 44156 42868 44158
rect 43820 44268 43876 44324
rect 41020 41468 41076 41524
rect 40684 37938 40740 37940
rect 40684 37886 40686 37938
rect 40686 37886 40738 37938
rect 40738 37886 40740 37938
rect 40684 37884 40740 37886
rect 41132 37826 41188 37828
rect 41132 37774 41134 37826
rect 41134 37774 41186 37826
rect 41186 37774 41188 37826
rect 41132 37772 41188 37774
rect 41244 36258 41300 36260
rect 41244 36206 41246 36258
rect 41246 36206 41298 36258
rect 41298 36206 41300 36258
rect 41244 36204 41300 36206
rect 41244 35980 41300 36036
rect 40684 34802 40740 34804
rect 40684 34750 40686 34802
rect 40686 34750 40738 34802
rect 40738 34750 40740 34802
rect 40684 34748 40740 34750
rect 41020 34748 41076 34804
rect 40124 33180 40180 33236
rect 39676 30098 39732 30100
rect 39676 30046 39678 30098
rect 39678 30046 39730 30098
rect 39730 30046 39732 30098
rect 39676 30044 39732 30046
rect 39564 28754 39620 28756
rect 39564 28702 39566 28754
rect 39566 28702 39618 28754
rect 39618 28702 39620 28754
rect 39564 28700 39620 28702
rect 39340 26012 39396 26068
rect 39340 25506 39396 25508
rect 39340 25454 39342 25506
rect 39342 25454 39394 25506
rect 39394 25454 39396 25506
rect 39340 25452 39396 25454
rect 40348 32732 40404 32788
rect 42140 34802 42196 34804
rect 42140 34750 42142 34802
rect 42142 34750 42194 34802
rect 42194 34750 42196 34802
rect 42140 34748 42196 34750
rect 41020 32284 41076 32340
rect 41132 31276 41188 31332
rect 40236 27858 40292 27860
rect 40236 27806 40238 27858
rect 40238 27806 40290 27858
rect 40290 27806 40292 27858
rect 40236 27804 40292 27806
rect 40236 26908 40292 26964
rect 39676 24668 39732 24724
rect 39788 24498 39844 24500
rect 39788 24446 39790 24498
rect 39790 24446 39842 24498
rect 39842 24446 39844 24498
rect 39788 24444 39844 24446
rect 40012 25564 40068 25620
rect 39676 20188 39732 20244
rect 40124 25506 40180 25508
rect 40124 25454 40126 25506
rect 40126 25454 40178 25506
rect 40178 25454 40180 25506
rect 40124 25452 40180 25454
rect 40124 23884 40180 23940
rect 39228 19852 39284 19908
rect 39228 18956 39284 19012
rect 39116 17388 39172 17444
rect 38668 15820 38724 15876
rect 39228 15820 39284 15876
rect 37436 4956 37492 5012
rect 40124 19906 40180 19908
rect 40124 19854 40126 19906
rect 40126 19854 40178 19906
rect 40178 19854 40180 19906
rect 40124 19852 40180 19854
rect 39900 17388 39956 17444
rect 39900 16044 39956 16100
rect 39788 4956 39844 5012
rect 40460 23938 40516 23940
rect 40460 23886 40462 23938
rect 40462 23886 40514 23938
rect 40514 23886 40516 23938
rect 40460 23884 40516 23886
rect 41692 31276 41748 31332
rect 41244 31218 41300 31220
rect 41244 31166 41246 31218
rect 41246 31166 41298 31218
rect 41298 31166 41300 31218
rect 41244 31164 41300 31166
rect 42364 31276 42420 31332
rect 41804 31164 41860 31220
rect 42588 31164 42644 31220
rect 44604 46114 44660 46116
rect 44604 46062 44606 46114
rect 44606 46062 44658 46114
rect 44658 46062 44660 46114
rect 44604 46060 44660 46062
rect 44828 45330 44884 45332
rect 44828 45278 44830 45330
rect 44830 45278 44882 45330
rect 44882 45278 44884 45330
rect 44828 45276 44884 45278
rect 44380 44492 44436 44548
rect 44828 44322 44884 44324
rect 44828 44270 44830 44322
rect 44830 44270 44882 44322
rect 44882 44270 44884 44322
rect 44828 44268 44884 44270
rect 44604 42812 44660 42868
rect 45612 43538 45668 43540
rect 45612 43486 45614 43538
rect 45614 43486 45666 43538
rect 45666 43486 45668 43538
rect 45612 43484 45668 43486
rect 45836 44546 45892 44548
rect 45836 44494 45838 44546
rect 45838 44494 45890 44546
rect 45890 44494 45892 44546
rect 45836 44492 45892 44494
rect 45724 43372 45780 43428
rect 46620 43426 46676 43428
rect 46620 43374 46622 43426
rect 46622 43374 46674 43426
rect 46674 43374 46676 43426
rect 46620 43372 46676 43374
rect 48188 46396 48244 46452
rect 47852 44380 47908 44436
rect 47628 41074 47684 41076
rect 47628 41022 47630 41074
rect 47630 41022 47682 41074
rect 47682 41022 47684 41074
rect 47628 41020 47684 41022
rect 48188 41074 48244 41076
rect 48188 41022 48190 41074
rect 48190 41022 48242 41074
rect 48242 41022 48244 41074
rect 48188 41020 48244 41022
rect 46172 38668 46228 38724
rect 43932 36204 43988 36260
rect 44492 37212 44548 37268
rect 43148 31052 43204 31108
rect 42028 30268 42084 30324
rect 41916 27804 41972 27860
rect 42028 25452 42084 25508
rect 43372 25340 43428 25396
rect 41244 24444 41300 24500
rect 41132 19292 41188 19348
rect 42028 4956 42084 5012
rect 40348 4562 40404 4564
rect 40348 4510 40350 4562
rect 40350 4510 40402 4562
rect 40402 4510 40404 4562
rect 40348 4508 40404 4510
rect 41244 4508 41300 4564
rect 41020 4060 41076 4116
rect 39004 3612 39060 3668
rect 40012 3666 40068 3668
rect 40012 3614 40014 3666
rect 40014 3614 40066 3666
rect 40066 3614 40068 3666
rect 40012 3612 40068 3614
rect 42252 4114 42308 4116
rect 42252 4062 42254 4114
rect 42254 4062 42306 4114
rect 42306 4062 42308 4114
rect 42252 4060 42308 4062
rect 42028 3612 42084 3668
rect 42812 3666 42868 3668
rect 42812 3614 42814 3666
rect 42814 3614 42866 3666
rect 42866 3614 42868 3666
rect 42812 3612 42868 3614
rect 44492 4508 44548 4564
rect 45052 25228 45108 25284
rect 43484 3500 43540 3556
rect 47852 37996 47908 38052
rect 47628 36370 47684 36372
rect 47628 36318 47630 36370
rect 47630 36318 47682 36370
rect 47682 36318 47684 36370
rect 47628 36316 47684 36318
rect 48188 36370 48244 36372
rect 48188 36318 48190 36370
rect 48190 36318 48242 36370
rect 48242 36318 48244 36370
rect 48188 36316 48244 36318
rect 47852 36258 47908 36260
rect 47852 36206 47854 36258
rect 47854 36206 47906 36258
rect 47906 36206 47908 36258
rect 47852 36204 47908 36206
rect 48188 35644 48244 35700
rect 47852 31106 47908 31108
rect 47852 31054 47854 31106
rect 47854 31054 47906 31106
rect 47906 31054 47908 31106
rect 47852 31052 47908 31054
rect 48188 30268 48244 30324
rect 47852 25452 47908 25508
rect 47628 25282 47684 25284
rect 47628 25230 47630 25282
rect 47630 25230 47682 25282
rect 47682 25230 47684 25282
rect 47628 25228 47684 25230
rect 48188 25228 48244 25284
rect 48188 24892 48244 24948
rect 46172 20076 46228 20132
rect 46284 21532 46340 21588
rect 47852 20130 47908 20132
rect 47852 20078 47854 20130
rect 47854 20078 47906 20130
rect 47906 20078 47908 20130
rect 47852 20076 47908 20078
rect 48188 19516 48244 19572
rect 47852 14306 47908 14308
rect 47852 14254 47854 14306
rect 47854 14254 47906 14306
rect 47906 14254 47908 14306
rect 47852 14252 47908 14254
rect 47628 14140 47684 14196
rect 48188 14140 48244 14196
rect 47852 9154 47908 9156
rect 47852 9102 47854 9154
rect 47854 9102 47906 9154
rect 47906 9102 47908 9154
rect 47852 9100 47908 9102
rect 47628 8764 47684 8820
rect 48188 8764 48244 8820
rect 47852 4562 47908 4564
rect 47852 4510 47854 4562
rect 47854 4510 47906 4562
rect 47906 4510 47908 4562
rect 47852 4508 47908 4510
rect 46284 3612 46340 3668
rect 45724 3554 45780 3556
rect 45724 3502 45726 3554
rect 45726 3502 45778 3554
rect 45778 3502 45780 3554
rect 45724 3500 45780 3502
rect 46620 3554 46676 3556
rect 46620 3502 46622 3554
rect 46622 3502 46674 3554
rect 46674 3502 46676 3554
rect 46620 3500 46676 3502
rect 47852 3666 47908 3668
rect 47852 3614 47854 3666
rect 47854 3614 47906 3666
rect 47906 3614 47908 3666
rect 47852 3612 47908 3614
rect 48188 3388 48244 3444
<< metal3 >>
rect 0 47572 800 47600
rect 0 47516 4844 47572
rect 4900 47516 4910 47572
rect 0 47488 800 47516
rect 2706 46844 2716 46900
rect 2772 46844 5628 46900
rect 5684 46844 5694 46900
rect 49200 46452 50000 46480
rect 48178 46396 48188 46452
rect 48244 46396 50000 46452
rect 49200 46368 50000 46396
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 28242 46060 28252 46116
rect 28308 46060 29484 46116
rect 29540 46060 29550 46116
rect 30930 46060 30940 46116
rect 30996 46060 33180 46116
rect 33236 46060 33246 46116
rect 33618 46060 33628 46116
rect 33684 46060 36988 46116
rect 37044 46060 37054 46116
rect 37650 46060 37660 46116
rect 37716 46060 40796 46116
rect 40852 46060 40862 46116
rect 41682 46060 41692 46116
rect 41748 46060 44604 46116
rect 44660 46060 44670 46116
rect 0 46004 800 46032
rect 0 45948 1932 46004
rect 1988 45948 1998 46004
rect 5618 45948 5628 46004
rect 5684 45948 6636 46004
rect 6692 45948 6702 46004
rect 0 45920 800 45948
rect 4722 45836 4732 45892
rect 4788 45836 5404 45892
rect 5460 45836 5470 45892
rect 16370 45836 16380 45892
rect 16436 45836 17052 45892
rect 17108 45836 17118 45892
rect 24098 45836 24108 45892
rect 24164 45836 25228 45892
rect 25284 45836 25294 45892
rect 33058 45836 33068 45892
rect 33124 45836 35980 45892
rect 36036 45836 36046 45892
rect 18946 45724 18956 45780
rect 19012 45724 21756 45780
rect 21812 45724 21822 45780
rect 7186 45612 7196 45668
rect 7252 45612 8428 45668
rect 8484 45612 8494 45668
rect 15250 45612 15260 45668
rect 15316 45612 23100 45668
rect 23156 45612 23166 45668
rect 4274 45500 4284 45556
rect 4340 45500 11676 45556
rect 11732 45500 11742 45556
rect 38612 45500 39788 45556
rect 39844 45500 39854 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 38612 45444 38668 45500
rect 18274 45388 18284 45444
rect 18340 45388 19068 45444
rect 19124 45388 19134 45444
rect 30268 45388 38668 45444
rect 30268 45332 30324 45388
rect 26898 45276 26908 45332
rect 26964 45276 28140 45332
rect 28196 45276 28206 45332
rect 28466 45276 28476 45332
rect 28532 45276 30324 45332
rect 34962 45276 34972 45332
rect 35028 45276 36988 45332
rect 37044 45276 37054 45332
rect 40338 45276 40348 45332
rect 40404 45276 41916 45332
rect 41972 45276 41982 45332
rect 43026 45276 43036 45332
rect 43092 45276 44828 45332
rect 44884 45276 44894 45332
rect 7858 45164 7868 45220
rect 7924 45164 8428 45220
rect 8642 45164 8652 45220
rect 8708 45164 14700 45220
rect 14756 45164 14766 45220
rect 25890 45164 25900 45220
rect 25956 45164 26908 45220
rect 8372 45108 8428 45164
rect 26852 45108 26908 45164
rect 8372 45052 12236 45108
rect 12292 45052 12302 45108
rect 24322 45052 24332 45108
rect 24388 45052 25564 45108
rect 25620 45052 25630 45108
rect 26852 45052 27132 45108
rect 27188 45052 27198 45108
rect 34402 45052 34412 45108
rect 34468 45052 35196 45108
rect 35252 45052 35262 45108
rect 32274 44940 32284 44996
rect 32340 44940 33292 44996
rect 33348 44940 33358 44996
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 24210 44492 24220 44548
rect 24276 44492 25452 44548
rect 25508 44492 25518 44548
rect 29586 44492 29596 44548
rect 29652 44492 30828 44548
rect 30884 44492 30894 44548
rect 36306 44492 36316 44548
rect 36372 44492 37996 44548
rect 38052 44492 38062 44548
rect 38994 44492 39004 44548
rect 39060 44492 40908 44548
rect 40964 44492 40974 44548
rect 44370 44492 44380 44548
rect 44436 44492 45836 44548
rect 45892 44492 45902 44548
rect 0 44436 800 44464
rect 0 44380 1820 44436
rect 1876 44380 1886 44436
rect 2044 44380 8092 44436
rect 8148 44380 8158 44436
rect 27430 44380 27468 44436
rect 27524 44380 27916 44436
rect 27972 44380 27982 44436
rect 41570 44380 41580 44436
rect 41636 44380 47852 44436
rect 47908 44380 47918 44436
rect 0 44352 800 44380
rect 2044 44324 2100 44380
rect 1586 44268 1596 44324
rect 1652 44268 2100 44324
rect 4834 44268 4844 44324
rect 4900 44268 5628 44324
rect 5684 44268 5964 44324
rect 6020 44268 6030 44324
rect 6188 44268 11340 44324
rect 11396 44268 11406 44324
rect 22754 44268 22764 44324
rect 22820 44268 24444 44324
rect 24500 44268 24510 44324
rect 35634 44268 35644 44324
rect 35700 44268 36988 44324
rect 37044 44268 37054 44324
rect 43810 44268 43820 44324
rect 43876 44268 44828 44324
rect 44884 44268 44894 44324
rect 6188 44100 6244 44268
rect 20962 44156 20972 44212
rect 21028 44156 22428 44212
rect 22484 44156 22494 44212
rect 30594 44156 30604 44212
rect 30660 44156 33404 44212
rect 33460 44156 33470 44212
rect 33730 44156 33740 44212
rect 33796 44156 39900 44212
rect 39956 44156 39966 44212
rect 41906 44156 41916 44212
rect 41972 44156 42812 44212
rect 42868 44156 42878 44212
rect 4274 44044 4284 44100
rect 4340 44044 6244 44100
rect 8372 44044 14812 44100
rect 14868 44044 14878 44100
rect 8372 43988 8428 44044
rect 4946 43932 4956 43988
rect 5012 43932 7420 43988
rect 7476 43932 7486 43988
rect 8082 43932 8092 43988
rect 8148 43932 8428 43988
rect 15092 43876 15148 44100
rect 15204 44044 15214 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 1474 43820 1484 43876
rect 1540 43820 15148 43876
rect 5618 43708 5628 43764
rect 5684 43708 6132 43764
rect 33394 43708 33404 43764
rect 33460 43708 35980 43764
rect 36036 43708 36046 43764
rect 6076 43652 6132 43708
rect 6076 43596 9324 43652
rect 9380 43596 9390 43652
rect 10546 43596 10556 43652
rect 10612 43596 12012 43652
rect 12068 43596 14252 43652
rect 14308 43596 14318 43652
rect 16370 43596 16380 43652
rect 16436 43596 17948 43652
rect 18004 43596 18014 43652
rect 18498 43596 18508 43652
rect 18564 43596 19180 43652
rect 19236 43596 21308 43652
rect 21364 43596 21868 43652
rect 21924 43596 21934 43652
rect 31602 43596 31612 43652
rect 31668 43596 38668 43652
rect 9426 43372 9436 43428
rect 9492 43372 11340 43428
rect 11396 43372 14812 43428
rect 14868 43372 14878 43428
rect 17948 43204 18004 43596
rect 38612 43540 38668 43596
rect 29586 43484 29596 43540
rect 29652 43484 31276 43540
rect 31332 43484 31342 43540
rect 33170 43484 33180 43540
rect 33236 43484 37324 43540
rect 37380 43484 37390 43540
rect 38612 43484 45612 43540
rect 45668 43484 45678 43540
rect 20402 43372 20412 43428
rect 20468 43372 21532 43428
rect 21588 43372 21598 43428
rect 28242 43372 28252 43428
rect 28308 43372 29036 43428
rect 29092 43372 29932 43428
rect 29988 43372 29998 43428
rect 45714 43372 45724 43428
rect 45780 43372 46620 43428
rect 46676 43372 46686 43428
rect 18162 43260 18172 43316
rect 18228 43260 18732 43316
rect 18788 43260 19404 43316
rect 19460 43260 19470 43316
rect 17948 43148 20636 43204
rect 20692 43148 20702 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 11106 43036 11116 43092
rect 11172 43036 21420 43092
rect 21476 43036 21868 43092
rect 21924 43036 23996 43092
rect 24052 43036 24780 43092
rect 24836 43036 24846 43092
rect 18022 42924 18060 42980
rect 18116 42924 18126 42980
rect 28914 42924 28924 42980
rect 28980 42924 29372 42980
rect 29428 42924 29438 42980
rect 0 42868 800 42896
rect 0 42812 1932 42868
rect 1988 42812 1998 42868
rect 2146 42812 2156 42868
rect 2212 42812 7028 42868
rect 8082 42812 8092 42868
rect 8148 42812 8988 42868
rect 9044 42812 9054 42868
rect 11554 42812 11564 42868
rect 11620 42812 12684 42868
rect 12740 42812 12750 42868
rect 17266 42812 17276 42868
rect 17332 42812 17342 42868
rect 19730 42812 19740 42868
rect 19796 42812 44604 42868
rect 44660 42812 44670 42868
rect 0 42784 800 42812
rect 6972 42756 7028 42812
rect 17276 42756 17332 42812
rect 4274 42700 4284 42756
rect 4340 42700 6748 42756
rect 6804 42700 6814 42756
rect 6972 42700 8148 42756
rect 8754 42700 8764 42756
rect 8820 42700 9996 42756
rect 10052 42700 10062 42756
rect 17276 42700 28476 42756
rect 28532 42700 29260 42756
rect 29316 42700 29326 42756
rect 8092 42644 8148 42700
rect 3938 42588 3948 42644
rect 4004 42588 7756 42644
rect 7812 42588 7822 42644
rect 8082 42588 8092 42644
rect 8148 42588 8158 42644
rect 7634 42476 7644 42532
rect 7700 42476 8428 42532
rect 8484 42476 8494 42532
rect 8764 42420 8820 42700
rect 9538 42588 9548 42644
rect 9604 42588 9884 42644
rect 9940 42588 13580 42644
rect 13636 42588 16604 42644
rect 16660 42588 17836 42644
rect 17892 42588 18508 42644
rect 18564 42588 18574 42644
rect 39778 42588 39788 42644
rect 39844 42588 40796 42644
rect 40852 42588 40862 42644
rect 8978 42476 8988 42532
rect 9044 42476 9660 42532
rect 9716 42476 9726 42532
rect 15474 42476 15484 42532
rect 15540 42476 16380 42532
rect 16436 42476 16446 42532
rect 18050 42476 18060 42532
rect 18116 42476 18396 42532
rect 18452 42476 18462 42532
rect 19506 42476 19516 42532
rect 19572 42476 23884 42532
rect 23940 42476 23950 42532
rect 29026 42476 29036 42532
rect 29092 42476 29260 42532
rect 29316 42476 29326 42532
rect 39218 42476 39228 42532
rect 39284 42476 40236 42532
rect 40292 42476 40908 42532
rect 40964 42476 40974 42532
rect 8082 42364 8092 42420
rect 8148 42364 8820 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 17388 42252 18844 42308
rect 18900 42252 19404 42308
rect 19460 42252 19470 42308
rect 22418 42252 22428 42308
rect 22484 42252 26908 42308
rect 17388 42196 17444 42252
rect 16930 42140 16940 42196
rect 16996 42140 17388 42196
rect 17444 42140 17454 42196
rect 18498 42140 18508 42196
rect 18564 42140 20076 42196
rect 20132 42140 21756 42196
rect 21812 42140 22204 42196
rect 22260 42140 22270 42196
rect 22642 42140 22652 42196
rect 22708 42140 22718 42196
rect 23426 42140 23436 42196
rect 23492 42140 26012 42196
rect 26068 42140 26078 42196
rect 8418 42028 8428 42084
rect 8484 42028 9324 42084
rect 9380 42028 9390 42084
rect 9986 42028 9996 42084
rect 10052 42028 11452 42084
rect 11508 42028 11518 42084
rect 14690 42028 14700 42084
rect 14756 42028 15036 42084
rect 15092 42028 18396 42084
rect 18452 42028 18462 42084
rect 18834 42028 18844 42084
rect 18900 42028 19516 42084
rect 19572 42028 19582 42084
rect 7298 41916 7308 41972
rect 7364 41916 8652 41972
rect 8708 41916 8718 41972
rect 10658 41916 10668 41972
rect 10724 41916 11900 41972
rect 11956 41916 11966 41972
rect 19394 41916 19404 41972
rect 19460 41916 20748 41972
rect 20804 41916 20814 41972
rect 22652 41860 22708 42140
rect 26852 42084 26908 42252
rect 26852 42028 27692 42084
rect 27748 42028 28140 42084
rect 28196 42028 28206 42084
rect 25330 41916 25340 41972
rect 25396 41916 27916 41972
rect 27972 41916 28476 41972
rect 28532 41916 28542 41972
rect 4498 41804 4508 41860
rect 4564 41804 7420 41860
rect 7476 41804 7486 41860
rect 8194 41804 8204 41860
rect 8260 41804 13580 41860
rect 13636 41804 13646 41860
rect 18386 41804 18396 41860
rect 18452 41804 18732 41860
rect 18788 41804 18798 41860
rect 22652 41804 23884 41860
rect 23940 41804 27580 41860
rect 27636 41804 27646 41860
rect 31154 41804 31164 41860
rect 31220 41804 32508 41860
rect 32564 41804 32574 41860
rect 10882 41692 10892 41748
rect 10948 41692 11340 41748
rect 11396 41692 11406 41748
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 11666 41468 11676 41524
rect 11732 41468 12460 41524
rect 12516 41468 12526 41524
rect 39778 41468 39788 41524
rect 39844 41468 41020 41524
rect 41076 41468 41086 41524
rect 2034 41356 2044 41412
rect 2100 41356 2110 41412
rect 10770 41356 10780 41412
rect 10836 41356 11900 41412
rect 11956 41356 11966 41412
rect 12684 41356 15148 41412
rect 22866 41356 22876 41412
rect 22932 41356 23548 41412
rect 23604 41356 23614 41412
rect 30482 41356 30492 41412
rect 30548 41356 32732 41412
rect 32788 41356 32798 41412
rect 0 41300 800 41328
rect 2044 41300 2100 41356
rect 12684 41300 12740 41356
rect 0 41244 2100 41300
rect 4834 41244 4844 41300
rect 4900 41244 5516 41300
rect 5572 41244 6972 41300
rect 7028 41244 7038 41300
rect 8866 41244 8876 41300
rect 8932 41244 9212 41300
rect 9268 41244 12740 41300
rect 15092 41300 15148 41356
rect 15092 41244 22988 41300
rect 23044 41244 23772 41300
rect 23828 41244 23838 41300
rect 0 41216 800 41244
rect 8978 41132 8988 41188
rect 9044 41132 12012 41188
rect 12068 41132 12572 41188
rect 12628 41132 13020 41188
rect 13076 41132 13086 41188
rect 18498 41132 18508 41188
rect 18564 41132 26124 41188
rect 26180 41132 26190 41188
rect 27570 41132 27580 41188
rect 27636 41132 28476 41188
rect 28532 41132 28542 41188
rect 49200 41076 50000 41104
rect 11890 41020 11900 41076
rect 11956 41020 15148 41076
rect 18162 41020 18172 41076
rect 18228 41020 18732 41076
rect 18788 41020 20412 41076
rect 20468 41020 22540 41076
rect 22596 41020 23100 41076
rect 23156 41020 23166 41076
rect 47618 41020 47628 41076
rect 47684 41020 48188 41076
rect 48244 41020 50000 41076
rect 15092 40964 15148 41020
rect 49200 40992 50000 41020
rect 2034 40908 2044 40964
rect 2100 40908 3836 40964
rect 3892 40908 5628 40964
rect 5684 40908 6860 40964
rect 6916 40908 6926 40964
rect 15092 40908 22148 40964
rect 22306 40908 22316 40964
rect 22372 40908 22652 40964
rect 22708 40908 25228 40964
rect 25284 40908 25294 40964
rect 27122 40908 27132 40964
rect 27188 40908 28140 40964
rect 28196 40908 28588 40964
rect 28644 40908 30716 40964
rect 30772 40908 30782 40964
rect 13794 40796 13804 40852
rect 13860 40796 14364 40852
rect 14420 40796 18900 40852
rect 8418 40684 8428 40740
rect 8484 40684 8494 40740
rect 8978 40684 8988 40740
rect 9044 40684 17724 40740
rect 17780 40684 18620 40740
rect 18676 40684 18686 40740
rect 8428 40516 8484 40684
rect 18844 40628 18900 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 22092 40740 22148 40908
rect 22092 40684 26572 40740
rect 26628 40684 27580 40740
rect 27636 40684 27646 40740
rect 12450 40572 12460 40628
rect 12516 40572 13692 40628
rect 13748 40572 18508 40628
rect 18564 40572 18574 40628
rect 18844 40572 22092 40628
rect 22148 40572 22158 40628
rect 27020 40572 29148 40628
rect 29204 40572 29214 40628
rect 27020 40516 27076 40572
rect 6626 40460 6636 40516
rect 6692 40460 7084 40516
rect 7140 40460 10668 40516
rect 10724 40460 10734 40516
rect 16818 40460 16828 40516
rect 16884 40460 27020 40516
rect 27076 40460 27086 40516
rect 8418 40348 8428 40404
rect 8484 40348 8988 40404
rect 9044 40348 9054 40404
rect 13346 40348 13356 40404
rect 13412 40348 13916 40404
rect 13972 40348 16380 40404
rect 16436 40348 16446 40404
rect 18050 40348 18060 40404
rect 18116 40348 19292 40404
rect 19348 40348 25004 40404
rect 25060 40348 25070 40404
rect 27570 40348 27580 40404
rect 27636 40348 28588 40404
rect 28644 40348 28654 40404
rect 4274 40236 4284 40292
rect 4340 40236 6748 40292
rect 6804 40236 6814 40292
rect 26898 40236 26908 40292
rect 26964 40236 28028 40292
rect 28084 40236 28094 40292
rect 31714 40236 31724 40292
rect 31780 40236 34188 40292
rect 34244 40236 34254 40292
rect 30706 40124 30716 40180
rect 30772 40124 31500 40180
rect 31556 40124 31566 40180
rect 29138 40012 29148 40068
rect 29204 40012 35028 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 7186 39900 7196 39956
rect 7252 39900 8204 39956
rect 8260 39900 8270 39956
rect 13906 39900 13916 39956
rect 13972 39900 30828 39956
rect 30884 39900 30894 39956
rect 34972 39844 35028 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 26852 39788 27132 39844
rect 27188 39788 27198 39844
rect 27458 39788 27468 39844
rect 27524 39788 27534 39844
rect 27906 39788 27916 39844
rect 27972 39788 27982 39844
rect 28802 39788 28812 39844
rect 28868 39788 32284 39844
rect 32340 39788 32350 39844
rect 34934 39788 34972 39844
rect 35028 39788 35532 39844
rect 35588 39788 35598 39844
rect 0 39732 800 39760
rect 26852 39732 26908 39788
rect 0 39676 1932 39732
rect 1988 39676 1998 39732
rect 15026 39676 15036 39732
rect 15092 39676 15708 39732
rect 15764 39676 15774 39732
rect 16034 39676 16044 39732
rect 16100 39676 16828 39732
rect 16884 39676 16894 39732
rect 20972 39676 26908 39732
rect 0 39648 800 39676
rect 20972 39620 21028 39676
rect 7298 39564 7308 39620
rect 7364 39564 10220 39620
rect 10276 39564 10892 39620
rect 10948 39564 10958 39620
rect 13682 39564 13692 39620
rect 13748 39564 21028 39620
rect 22306 39564 22316 39620
rect 22372 39564 23212 39620
rect 23268 39564 26908 39620
rect 26964 39564 26974 39620
rect 5282 39452 5292 39508
rect 5348 39452 6748 39508
rect 6804 39452 6814 39508
rect 20290 39452 20300 39508
rect 20356 39452 21980 39508
rect 22036 39452 22046 39508
rect 22754 39452 22764 39508
rect 22820 39452 23772 39508
rect 23828 39452 23838 39508
rect 27468 39396 27524 39788
rect 27916 39620 27972 39788
rect 28130 39676 28140 39732
rect 28196 39676 30156 39732
rect 30212 39676 30222 39732
rect 27916 39564 29484 39620
rect 29540 39564 32732 39620
rect 32788 39564 35980 39620
rect 36036 39564 36046 39620
rect 14130 39340 14140 39396
rect 14196 39340 16156 39396
rect 16212 39340 16716 39396
rect 16772 39340 16782 39396
rect 19618 39340 19628 39396
rect 19684 39340 20636 39396
rect 20692 39340 21308 39396
rect 21364 39340 21374 39396
rect 21634 39340 21644 39396
rect 21700 39340 22428 39396
rect 22484 39340 26460 39396
rect 26516 39340 26908 39396
rect 26964 39340 27524 39396
rect 14242 39228 14252 39284
rect 14308 39228 15148 39284
rect 27346 39228 27356 39284
rect 27412 39228 28812 39284
rect 28868 39228 28878 39284
rect 15092 39172 15148 39228
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 14354 39116 14364 39172
rect 14420 39116 14700 39172
rect 14756 39116 14766 39172
rect 15092 39116 16268 39172
rect 16324 39116 18060 39172
rect 18116 39116 18126 39172
rect 27570 39116 27580 39172
rect 27636 39116 33404 39172
rect 33460 39116 33470 39172
rect 8530 39004 8540 39060
rect 8596 39004 9436 39060
rect 9492 39004 9502 39060
rect 12562 39004 12572 39060
rect 12628 39004 13916 39060
rect 13972 39004 13982 39060
rect 16482 39004 16492 39060
rect 16548 39004 17388 39060
rect 17444 39004 27188 39060
rect 27346 39004 27356 39060
rect 27412 39004 28252 39060
rect 28308 39004 28318 39060
rect 28690 39004 28700 39060
rect 28756 39004 29372 39060
rect 29428 39004 29438 39060
rect 30818 39004 30828 39060
rect 30884 39004 32508 39060
rect 32564 39004 32574 39060
rect 27132 38948 27188 39004
rect 12450 38892 12460 38948
rect 12516 38892 13468 38948
rect 13524 38892 13534 38948
rect 18834 38892 18844 38948
rect 18900 38892 20300 38948
rect 20356 38892 20366 38948
rect 23986 38892 23996 38948
rect 24052 38892 26908 38948
rect 27132 38892 34524 38948
rect 34580 38892 36092 38948
rect 36148 38892 36158 38948
rect 26852 38836 26908 38892
rect 9874 38780 9884 38836
rect 9940 38780 10556 38836
rect 10612 38780 11676 38836
rect 11732 38780 11742 38836
rect 12114 38780 12124 38836
rect 12180 38780 13692 38836
rect 13748 38780 13758 38836
rect 14578 38780 14588 38836
rect 14644 38780 15036 38836
rect 15092 38780 17836 38836
rect 17892 38780 18620 38836
rect 18676 38780 18686 38836
rect 24658 38780 24668 38836
rect 24724 38780 25340 38836
rect 25396 38780 25406 38836
rect 26852 38780 27916 38836
rect 27972 38780 29204 38836
rect 3826 38668 3836 38724
rect 3892 38668 4844 38724
rect 4900 38668 4910 38724
rect 11890 38668 11900 38724
rect 11956 38668 14700 38724
rect 14756 38668 14766 38724
rect 18498 38668 18508 38724
rect 18564 38668 19180 38724
rect 19236 38668 19246 38724
rect 26562 38668 26572 38724
rect 26628 38668 27020 38724
rect 27076 38668 28252 38724
rect 28308 38668 28318 38724
rect 12460 38556 17052 38612
rect 17108 38556 17118 38612
rect 27346 38556 27356 38612
rect 27412 38556 27468 38612
rect 27524 38556 27534 38612
rect 27682 38556 27692 38612
rect 27748 38556 27916 38612
rect 27972 38556 27982 38612
rect 12460 38500 12516 38556
rect 29148 38500 29204 38780
rect 30706 38668 30716 38724
rect 30772 38668 33292 38724
rect 33348 38668 33358 38724
rect 34290 38668 34300 38724
rect 34356 38668 36652 38724
rect 36708 38668 46172 38724
rect 46228 38668 46238 38724
rect 11890 38444 11900 38500
rect 11956 38444 12460 38500
rect 12516 38444 12526 38500
rect 26786 38444 26796 38500
rect 26852 38444 27692 38500
rect 27748 38444 27758 38500
rect 29138 38444 29148 38500
rect 29204 38444 29214 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 14354 38332 14364 38388
rect 14420 38332 17612 38388
rect 17668 38332 17678 38388
rect 2828 38220 9996 38276
rect 10052 38220 10062 38276
rect 0 38164 800 38192
rect 2828 38164 2884 38220
rect 0 38108 1932 38164
rect 1988 38108 1998 38164
rect 2146 38108 2156 38164
rect 2212 38108 2828 38164
rect 2884 38108 2894 38164
rect 4918 38108 4956 38164
rect 5012 38108 5022 38164
rect 10434 38108 10444 38164
rect 10500 38108 11116 38164
rect 11172 38108 19404 38164
rect 19460 38108 19470 38164
rect 0 38080 800 38108
rect 3266 37996 3276 38052
rect 3332 37940 3388 38052
rect 4274 37996 4284 38052
rect 4340 37996 7644 38052
rect 7700 37996 7710 38052
rect 13906 37996 13916 38052
rect 13972 37996 27132 38052
rect 27188 37996 27198 38052
rect 39778 37996 39788 38052
rect 39844 37996 47852 38052
rect 47908 37996 47918 38052
rect 3332 37884 4844 37940
rect 4900 37884 4910 37940
rect 39106 37884 39116 37940
rect 39172 37884 39340 37940
rect 39396 37884 40684 37940
rect 40740 37884 40750 37940
rect 18722 37772 18732 37828
rect 18788 37772 20300 37828
rect 20356 37772 20366 37828
rect 21746 37772 21756 37828
rect 21812 37772 23212 37828
rect 23268 37772 23278 37828
rect 38994 37772 39004 37828
rect 39060 37772 41132 37828
rect 41188 37772 41198 37828
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 3602 37548 3612 37604
rect 3668 37548 4844 37604
rect 4900 37548 4910 37604
rect 5170 37436 5180 37492
rect 5236 37436 8092 37492
rect 8148 37436 13804 37492
rect 13860 37436 13870 37492
rect 27906 37436 27916 37492
rect 27972 37436 29372 37492
rect 29428 37436 29438 37492
rect 32498 37436 32508 37492
rect 32564 37436 33180 37492
rect 33236 37436 33246 37492
rect 9538 37324 9548 37380
rect 9604 37324 9996 37380
rect 10052 37324 12460 37380
rect 12516 37324 12796 37380
rect 12852 37324 13916 37380
rect 13972 37324 13982 37380
rect 18050 37324 18060 37380
rect 18116 37324 20524 37380
rect 20580 37324 20590 37380
rect 33730 37324 33740 37380
rect 33796 37324 34860 37380
rect 34916 37324 34926 37380
rect 2370 37212 2380 37268
rect 2436 37212 5628 37268
rect 5684 37212 5694 37268
rect 9548 37212 10220 37268
rect 10276 37212 10892 37268
rect 10948 37212 10958 37268
rect 12002 37212 12012 37268
rect 12068 37212 12572 37268
rect 12628 37212 12638 37268
rect 15810 37212 15820 37268
rect 15876 37212 21420 37268
rect 21476 37212 21486 37268
rect 28466 37212 28476 37268
rect 28532 37212 29932 37268
rect 29988 37212 44492 37268
rect 44548 37212 44558 37268
rect 9548 37156 9604 37212
rect 4274 37100 4284 37156
rect 4340 37100 7756 37156
rect 7812 37100 7822 37156
rect 8866 37100 8876 37156
rect 8932 37100 9548 37156
rect 9604 37100 9614 37156
rect 9762 37100 9772 37156
rect 9828 37100 9866 37156
rect 12674 37100 12684 37156
rect 12740 37100 13244 37156
rect 13300 37100 15148 37156
rect 15204 37100 15214 37156
rect 18834 37100 18844 37156
rect 18900 37100 19068 37156
rect 19124 37100 19134 37156
rect 33954 37100 33964 37156
rect 34020 37100 35420 37156
rect 35476 37100 35868 37156
rect 35924 37100 35934 37156
rect 4498 36988 4508 37044
rect 4564 36988 5180 37044
rect 5236 36988 8092 37044
rect 8148 36988 12460 37044
rect 12516 36988 12526 37044
rect 18498 36988 18508 37044
rect 18564 36988 19292 37044
rect 19348 36988 20076 37044
rect 20132 36988 20142 37044
rect 23538 36988 23548 37044
rect 23604 36988 33740 37044
rect 33796 36988 33806 37044
rect 4946 36876 4956 36932
rect 5012 36876 10500 36932
rect 10658 36876 10668 36932
rect 10724 36876 11452 36932
rect 11508 36876 11518 36932
rect 14018 36876 14028 36932
rect 14084 36876 14812 36932
rect 14868 36876 14878 36932
rect 16594 36876 16604 36932
rect 16660 36876 20300 36932
rect 20356 36876 27244 36932
rect 27300 36876 28140 36932
rect 28196 36876 28206 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 10444 36820 10500 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 4834 36764 4844 36820
rect 4900 36764 5628 36820
rect 5684 36764 5694 36820
rect 10444 36764 11564 36820
rect 11620 36764 11630 36820
rect 2930 36652 2940 36708
rect 2996 36652 5852 36708
rect 5908 36652 5918 36708
rect 12002 36652 12012 36708
rect 12068 36652 13356 36708
rect 13412 36652 13422 36708
rect 0 36596 800 36624
rect 0 36540 1932 36596
rect 1988 36540 1998 36596
rect 4050 36540 4060 36596
rect 4116 36540 5740 36596
rect 5796 36540 5806 36596
rect 11106 36540 11116 36596
rect 11172 36540 12236 36596
rect 12292 36540 12302 36596
rect 13122 36540 13132 36596
rect 13188 36540 13580 36596
rect 13636 36540 13646 36596
rect 13990 36540 14028 36596
rect 14084 36540 14094 36596
rect 15586 36540 15596 36596
rect 15652 36540 16156 36596
rect 16212 36540 16222 36596
rect 17154 36540 17164 36596
rect 17220 36540 20860 36596
rect 20916 36540 22652 36596
rect 22708 36540 22718 36596
rect 0 36512 800 36540
rect 4946 36428 4956 36484
rect 5012 36428 6076 36484
rect 6132 36428 6142 36484
rect 8306 36428 8316 36484
rect 8372 36428 9884 36484
rect 9940 36428 12908 36484
rect 12964 36428 12974 36484
rect 13458 36428 13468 36484
rect 13524 36428 14812 36484
rect 14868 36428 14878 36484
rect 15474 36428 15484 36484
rect 15540 36428 19292 36484
rect 19348 36428 19358 36484
rect 5058 36316 5068 36372
rect 5124 36316 5516 36372
rect 5572 36316 8428 36372
rect 8484 36316 8494 36372
rect 11778 36316 11788 36372
rect 11844 36316 12684 36372
rect 12740 36316 12750 36372
rect 13692 36316 19180 36372
rect 19236 36316 19246 36372
rect 21186 36316 21196 36372
rect 21252 36316 22316 36372
rect 22372 36316 22382 36372
rect 47618 36316 47628 36372
rect 47684 36316 48188 36372
rect 48244 36316 48254 36372
rect 10882 36204 10892 36260
rect 10948 36204 13468 36260
rect 13524 36204 13534 36260
rect 13692 36148 13748 36316
rect 13878 36204 13916 36260
rect 13972 36204 13982 36260
rect 14802 36204 14812 36260
rect 14868 36204 15484 36260
rect 15540 36204 15550 36260
rect 16034 36204 16044 36260
rect 16100 36204 17948 36260
rect 18004 36204 18014 36260
rect 18834 36204 18844 36260
rect 18900 36204 19852 36260
rect 19908 36204 19918 36260
rect 22530 36204 22540 36260
rect 22596 36204 32172 36260
rect 32228 36204 34748 36260
rect 34804 36204 34814 36260
rect 41234 36204 41244 36260
rect 41300 36204 43932 36260
rect 43988 36204 43998 36260
rect 47842 36204 47852 36260
rect 47908 36204 47918 36260
rect 11218 36092 11228 36148
rect 11284 36092 11676 36148
rect 11732 36092 11742 36148
rect 12198 36092 12236 36148
rect 12292 36092 12302 36148
rect 12450 36092 12460 36148
rect 12516 36092 13748 36148
rect 13804 36092 16380 36148
rect 16436 36092 18620 36148
rect 18676 36092 18686 36148
rect 13804 36036 13860 36092
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 47852 36036 47908 36204
rect 11554 35980 11564 36036
rect 11620 35980 13860 36036
rect 13916 35980 19684 36036
rect 41234 35980 41244 36036
rect 41300 35980 47908 36036
rect 3042 35868 3052 35924
rect 3108 35868 3500 35924
rect 3556 35868 3566 35924
rect 10322 35868 10332 35924
rect 10388 35868 11676 35924
rect 11732 35868 11742 35924
rect 13916 35812 13972 35980
rect 19628 35924 19684 35980
rect 14690 35868 14700 35924
rect 14756 35868 15036 35924
rect 15092 35868 15708 35924
rect 15764 35868 15774 35924
rect 19590 35868 19628 35924
rect 19684 35868 22204 35924
rect 22260 35868 22876 35924
rect 22932 35868 22942 35924
rect 6178 35756 6188 35812
rect 6244 35756 13972 35812
rect 18050 35756 18060 35812
rect 18116 35756 18844 35812
rect 18900 35756 18910 35812
rect 19282 35756 19292 35812
rect 19348 35756 19740 35812
rect 19796 35756 38668 35812
rect 38724 35756 39004 35812
rect 39060 35756 39070 35812
rect 49200 35700 50000 35728
rect 9874 35644 9884 35700
rect 9940 35644 10668 35700
rect 10724 35644 10734 35700
rect 14018 35644 14028 35700
rect 14084 35644 14364 35700
rect 14420 35644 23548 35700
rect 23604 35644 23614 35700
rect 48178 35644 48188 35700
rect 48244 35644 50000 35700
rect 49200 35616 50000 35644
rect 13346 35532 13356 35588
rect 13412 35532 18844 35588
rect 18900 35532 18910 35588
rect 21970 35532 21980 35588
rect 22036 35532 23324 35588
rect 23380 35532 23390 35588
rect 32498 35532 32508 35588
rect 32564 35532 33852 35588
rect 33908 35532 33918 35588
rect 35074 35532 35084 35588
rect 35140 35532 35980 35588
rect 36036 35532 36046 35588
rect 2034 35420 2044 35476
rect 2100 35420 17500 35476
rect 17556 35420 18284 35476
rect 18340 35420 18350 35476
rect 18610 35420 18620 35476
rect 18676 35420 19292 35476
rect 19348 35420 19358 35476
rect 35522 35420 35532 35476
rect 35588 35420 37212 35476
rect 37268 35420 37278 35476
rect 7298 35308 7308 35364
rect 7364 35308 8316 35364
rect 8372 35308 8382 35364
rect 12338 35308 12348 35364
rect 12404 35308 13132 35364
rect 13188 35308 13198 35364
rect 16818 35308 16828 35364
rect 16884 35308 17388 35364
rect 17444 35308 18060 35364
rect 18116 35308 18126 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 9650 35196 9660 35252
rect 9716 35196 15932 35252
rect 15988 35196 15998 35252
rect 26852 35196 30492 35252
rect 30548 35196 30558 35252
rect 26852 35140 26908 35196
rect 4274 35084 4284 35140
rect 4340 35084 7308 35140
rect 7364 35084 7374 35140
rect 9762 35084 9772 35140
rect 9828 35084 10780 35140
rect 10836 35084 10846 35140
rect 12114 35084 12124 35140
rect 12180 35084 14028 35140
rect 14084 35084 14094 35140
rect 24882 35084 24892 35140
rect 24948 35084 26908 35140
rect 28578 35084 28588 35140
rect 28644 35084 30044 35140
rect 30100 35084 30828 35140
rect 30884 35084 30894 35140
rect 34514 35084 34524 35140
rect 34580 35084 39340 35140
rect 39396 35084 39406 35140
rect 0 35028 800 35056
rect 0 34972 1932 35028
rect 1988 34972 1998 35028
rect 3154 34972 3164 35028
rect 3220 34972 6468 35028
rect 6626 34972 6636 35028
rect 6692 34972 8540 35028
rect 8596 34972 13692 35028
rect 13748 34972 13758 35028
rect 0 34944 800 34972
rect 6412 34916 6468 34972
rect 2818 34860 2828 34916
rect 2884 34860 3612 34916
rect 3668 34860 3678 34916
rect 6412 34860 13468 34916
rect 13524 34860 13534 34916
rect 15092 34860 21644 34916
rect 21700 34860 22428 34916
rect 22484 34860 22876 34916
rect 22932 34860 22942 34916
rect 15092 34804 15148 34860
rect 2930 34748 2940 34804
rect 2996 34748 4396 34804
rect 4452 34748 4844 34804
rect 4900 34748 5628 34804
rect 5684 34748 5694 34804
rect 5954 34748 5964 34804
rect 6020 34748 7980 34804
rect 8036 34748 8046 34804
rect 9426 34748 9436 34804
rect 9492 34748 12572 34804
rect 12628 34748 12638 34804
rect 12898 34748 12908 34804
rect 12964 34748 15148 34804
rect 22306 34748 22316 34804
rect 22372 34748 23212 34804
rect 23268 34748 24556 34804
rect 24612 34748 24622 34804
rect 28588 34692 28644 35084
rect 29810 34972 29820 35028
rect 29876 34972 30268 35028
rect 30324 34972 30334 35028
rect 32722 34972 32732 35028
rect 32788 34972 36092 35028
rect 36148 34972 36158 35028
rect 29138 34748 29148 34804
rect 29204 34748 29708 34804
rect 29764 34748 30268 34804
rect 30324 34748 30334 34804
rect 40674 34748 40684 34804
rect 40740 34748 41020 34804
rect 41076 34748 42140 34804
rect 42196 34748 42206 34804
rect 18722 34636 18732 34692
rect 18788 34636 19180 34692
rect 19236 34636 23324 34692
rect 23380 34636 28644 34692
rect 11778 34524 11788 34580
rect 11844 34524 12236 34580
rect 12292 34524 12302 34580
rect 14466 34524 14476 34580
rect 14532 34524 15372 34580
rect 15428 34524 15438 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 20972 34412 28588 34468
rect 28644 34412 29820 34468
rect 29876 34412 29886 34468
rect 20972 34356 21028 34412
rect 12674 34300 12684 34356
rect 12740 34300 13132 34356
rect 13188 34300 21028 34356
rect 24434 34300 24444 34356
rect 24500 34300 25340 34356
rect 25396 34300 25406 34356
rect 2706 34188 2716 34244
rect 2772 34188 3052 34244
rect 3108 34188 26124 34244
rect 26180 34188 26190 34244
rect 16706 34076 16716 34132
rect 16772 34076 18284 34132
rect 18340 34076 18350 34132
rect 24994 34076 25004 34132
rect 25060 34076 26796 34132
rect 26852 34076 26908 34132
rect 26964 34076 26974 34132
rect 3602 33964 3612 34020
rect 3668 33964 4508 34020
rect 4564 33964 7644 34020
rect 7700 33964 7710 34020
rect 18498 33964 18508 34020
rect 18564 33964 19964 34020
rect 20020 33964 26124 34020
rect 26180 33964 26190 34020
rect 28242 33964 28252 34020
rect 28308 33964 33516 34020
rect 33572 33964 33582 34020
rect 29484 33852 35532 33908
rect 35588 33852 35598 33908
rect 29484 33796 29540 33852
rect 6402 33740 6412 33796
rect 6468 33740 7420 33796
rect 7476 33740 7486 33796
rect 29474 33740 29484 33796
rect 29540 33740 29550 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 21970 33628 21980 33684
rect 22036 33628 23100 33684
rect 23156 33628 24332 33684
rect 24388 33628 24398 33684
rect 28466 33628 28476 33684
rect 28532 33628 28542 33684
rect 28476 33572 28532 33628
rect 28476 33516 29148 33572
rect 29204 33516 29214 33572
rect 0 33460 800 33488
rect 0 33404 1708 33460
rect 1764 33404 2492 33460
rect 2548 33404 2558 33460
rect 12002 33404 12012 33460
rect 12068 33404 17724 33460
rect 17780 33404 17790 33460
rect 22838 33404 22876 33460
rect 22932 33404 22942 33460
rect 25218 33404 25228 33460
rect 25284 33404 26236 33460
rect 26292 33404 27020 33460
rect 27076 33404 27086 33460
rect 27570 33404 27580 33460
rect 27636 33404 28028 33460
rect 28084 33404 28588 33460
rect 28644 33404 28654 33460
rect 35522 33404 35532 33460
rect 35588 33404 38892 33460
rect 38948 33404 38958 33460
rect 0 33376 800 33404
rect 7970 33292 7980 33348
rect 8036 33292 9548 33348
rect 9604 33292 9614 33348
rect 9762 33292 9772 33348
rect 9828 33292 9996 33348
rect 10052 33292 10108 33348
rect 10164 33292 10174 33348
rect 12786 33292 12796 33348
rect 12852 33292 17668 33348
rect 17826 33292 17836 33348
rect 17892 33292 18508 33348
rect 18564 33292 26908 33348
rect 27682 33292 27692 33348
rect 27748 33292 29372 33348
rect 29428 33292 29438 33348
rect 30380 33292 35868 33348
rect 35924 33292 35934 33348
rect 17612 33236 17668 33292
rect 9762 33180 9772 33236
rect 9828 33180 17052 33236
rect 17108 33180 17118 33236
rect 17612 33180 18956 33236
rect 19012 33180 19022 33236
rect 22642 33180 22652 33236
rect 22708 33180 22988 33236
rect 23044 33180 23054 33236
rect 26852 33124 26908 33292
rect 30380 33236 30436 33292
rect 28242 33180 28252 33236
rect 28308 33180 29036 33236
rect 29092 33180 29102 33236
rect 29698 33180 29708 33236
rect 29764 33180 30380 33236
rect 30436 33180 30446 33236
rect 34066 33180 34076 33236
rect 34132 33180 35756 33236
rect 35812 33180 35822 33236
rect 38612 33180 40124 33236
rect 40180 33180 40190 33236
rect 38612 33124 38668 33180
rect 9874 33068 9884 33124
rect 9940 33068 10444 33124
rect 10500 33068 10510 33124
rect 26852 33068 38668 33124
rect 19394 32956 19404 33012
rect 19460 32956 19628 33012
rect 19684 32956 19694 33012
rect 34514 32956 34524 33012
rect 34580 32956 34860 33012
rect 34916 32956 34926 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 26898 32844 26908 32900
rect 26964 32844 27002 32900
rect 26786 32732 26796 32788
rect 10770 32620 10780 32676
rect 10836 32620 12348 32676
rect 12404 32620 12414 32676
rect 12674 32620 12684 32676
rect 12740 32620 13692 32676
rect 13748 32620 13758 32676
rect 26852 32620 26908 32788
rect 34374 32732 34412 32788
rect 34468 32732 34478 32788
rect 36866 32732 36876 32788
rect 36932 32732 40348 32788
rect 40404 32732 40414 32788
rect 26964 32620 26974 32676
rect 34514 32620 34524 32676
rect 34580 32620 34860 32676
rect 34916 32620 38668 32676
rect 10994 32508 11004 32564
rect 11060 32508 12460 32564
rect 12516 32508 12908 32564
rect 12964 32508 12974 32564
rect 14354 32508 14364 32564
rect 14420 32508 15596 32564
rect 15652 32508 17612 32564
rect 17668 32508 17678 32564
rect 35746 32508 35756 32564
rect 35812 32508 36428 32564
rect 36484 32508 36494 32564
rect 27010 32396 27020 32452
rect 27076 32396 28364 32452
rect 28420 32396 28430 32452
rect 36306 32396 36316 32452
rect 36372 32396 38220 32452
rect 38276 32396 38286 32452
rect 38612 32340 38668 32620
rect 9174 32284 9212 32340
rect 9268 32284 9278 32340
rect 10546 32284 10556 32340
rect 10612 32284 17612 32340
rect 17668 32284 17678 32340
rect 26852 32284 35420 32340
rect 35476 32284 36876 32340
rect 36932 32284 36942 32340
rect 38612 32284 41020 32340
rect 41076 32284 41086 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 10434 32060 10444 32116
rect 10500 32060 24444 32116
rect 24500 32060 24510 32116
rect 26852 32004 26908 32284
rect 28354 32172 28364 32228
rect 28420 32172 28700 32228
rect 28756 32172 28766 32228
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 27804 32060 29148 32116
rect 29204 32060 29708 32116
rect 29764 32060 29774 32116
rect 33842 32060 33852 32116
rect 33908 32060 34188 32116
rect 34244 32060 34254 32116
rect 27804 32004 27860 32060
rect 8194 31948 8204 32004
rect 8260 31948 9436 32004
rect 9492 31948 9884 32004
rect 9940 31948 10668 32004
rect 10724 31948 10734 32004
rect 23650 31948 23660 32004
rect 23716 31948 26908 32004
rect 27794 31948 27804 32004
rect 27860 31948 27870 32004
rect 33618 31948 33628 32004
rect 33684 31948 34748 32004
rect 34804 31948 36876 32004
rect 36932 31948 36942 32004
rect 0 31892 800 31920
rect 0 31836 1820 31892
rect 1876 31836 1886 31892
rect 5058 31836 5068 31892
rect 5124 31836 6636 31892
rect 6692 31836 6702 31892
rect 10098 31836 10108 31892
rect 10164 31836 10780 31892
rect 10836 31836 10846 31892
rect 13906 31836 13916 31892
rect 13972 31836 19404 31892
rect 19460 31836 19470 31892
rect 19842 31836 19852 31892
rect 19908 31836 21756 31892
rect 21812 31836 21822 31892
rect 23202 31836 23212 31892
rect 23268 31836 36988 31892
rect 37044 31836 37054 31892
rect 0 31808 800 31836
rect 1922 31724 1932 31780
rect 1988 31724 4284 31780
rect 4340 31724 5740 31780
rect 5796 31724 5806 31780
rect 9538 31724 9548 31780
rect 9604 31724 12124 31780
rect 12180 31724 12190 31780
rect 13346 31724 13356 31780
rect 13412 31724 14028 31780
rect 14084 31724 14094 31780
rect 18050 31724 18060 31780
rect 18116 31724 19068 31780
rect 19124 31724 19134 31780
rect 19292 31724 19740 31780
rect 19796 31724 19806 31780
rect 19954 31724 19964 31780
rect 20020 31724 27580 31780
rect 27636 31724 33852 31780
rect 33908 31724 33918 31780
rect 19292 31668 19348 31724
rect 4050 31612 4060 31668
rect 4116 31612 7980 31668
rect 8036 31612 8046 31668
rect 8316 31612 9324 31668
rect 9380 31612 9390 31668
rect 9650 31612 9660 31668
rect 9716 31612 13804 31668
rect 13860 31612 13870 31668
rect 18498 31612 18508 31668
rect 18564 31612 19348 31668
rect 25554 31612 25564 31668
rect 25620 31612 26908 31668
rect 27234 31612 27244 31668
rect 27300 31612 29036 31668
rect 29092 31612 29102 31668
rect 33618 31612 33628 31668
rect 33684 31612 34188 31668
rect 34244 31612 34254 31668
rect 8316 31556 8372 31612
rect 26852 31556 26908 31612
rect 5842 31500 5852 31556
rect 5908 31500 8092 31556
rect 8148 31500 8158 31556
rect 8306 31500 8316 31556
rect 8372 31500 8410 31556
rect 8530 31500 8540 31556
rect 8596 31500 8634 31556
rect 8866 31500 8876 31556
rect 8932 31500 9772 31556
rect 9828 31500 9838 31556
rect 12674 31500 12684 31556
rect 12740 31500 13468 31556
rect 13524 31500 13534 31556
rect 19058 31500 19068 31556
rect 19124 31500 23660 31556
rect 23716 31500 23726 31556
rect 26852 31500 27580 31556
rect 27636 31500 34076 31556
rect 34132 31500 34142 31556
rect 37090 31500 37100 31556
rect 37156 31500 37436 31556
rect 37492 31500 37502 31556
rect 7634 31388 7644 31444
rect 7700 31388 11228 31444
rect 11284 31388 11294 31444
rect 26898 31388 26908 31444
rect 26964 31388 27002 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 8726 31276 8764 31332
rect 8820 31276 8830 31332
rect 10210 31276 10220 31332
rect 10276 31276 16044 31332
rect 16100 31276 16110 31332
rect 20290 31276 20300 31332
rect 20356 31276 22764 31332
rect 22820 31276 41132 31332
rect 41188 31276 41692 31332
rect 41748 31276 42364 31332
rect 42420 31276 42430 31332
rect 6066 31164 6076 31220
rect 6132 31164 9436 31220
rect 9492 31164 9502 31220
rect 9874 31164 9884 31220
rect 9940 31164 11564 31220
rect 11620 31164 11630 31220
rect 14578 31164 14588 31220
rect 14644 31164 14654 31220
rect 19506 31164 19516 31220
rect 19572 31164 20412 31220
rect 20468 31164 20478 31220
rect 21522 31164 21532 31220
rect 21588 31164 23212 31220
rect 23268 31164 23278 31220
rect 32722 31164 32732 31220
rect 32788 31164 33740 31220
rect 33796 31164 34188 31220
rect 34244 31164 34254 31220
rect 36978 31164 36988 31220
rect 37044 31164 37996 31220
rect 38052 31164 41244 31220
rect 41300 31164 41804 31220
rect 41860 31164 42588 31220
rect 42644 31164 42654 31220
rect 14588 31108 14644 31164
rect 9090 31052 9100 31108
rect 9156 31052 11452 31108
rect 11508 31052 11518 31108
rect 14588 31052 15260 31108
rect 15316 31052 15326 31108
rect 18162 31052 18172 31108
rect 18228 31052 18844 31108
rect 18900 31052 19404 31108
rect 19460 31052 20300 31108
rect 20356 31052 20366 31108
rect 26852 31052 27356 31108
rect 27412 31052 30380 31108
rect 30436 31052 30446 31108
rect 33842 31052 33852 31108
rect 33908 31052 34860 31108
rect 34916 31052 34926 31108
rect 43138 31052 43148 31108
rect 43204 31052 47852 31108
rect 47908 31052 47918 31108
rect 7746 30940 7756 30996
rect 7812 30940 9772 30996
rect 9828 30940 9838 30996
rect 9986 30940 9996 30996
rect 10052 30940 10892 30996
rect 10948 30940 10958 30996
rect 11890 30940 11900 30996
rect 11956 30940 20636 30996
rect 20692 30940 20702 30996
rect 9996 30884 10052 30940
rect 3938 30828 3948 30884
rect 4004 30828 7644 30884
rect 7700 30828 7710 30884
rect 8530 30828 8540 30884
rect 8596 30828 10052 30884
rect 14214 30828 14252 30884
rect 14308 30828 14318 30884
rect 14466 30828 14476 30884
rect 14532 30828 17388 30884
rect 17444 30828 17454 30884
rect 8194 30716 8204 30772
rect 8260 30716 14812 30772
rect 14868 30716 14878 30772
rect 26852 30660 26908 31052
rect 28130 30940 28140 30996
rect 28196 30940 28588 30996
rect 28644 30940 28654 30996
rect 34066 30940 34076 30996
rect 34132 30940 36540 30996
rect 36596 30940 36606 30996
rect 34860 30884 34916 30940
rect 34850 30828 34860 30884
rect 34916 30828 34926 30884
rect 35970 30716 35980 30772
rect 36036 30716 36988 30772
rect 37044 30716 37054 30772
rect 19618 30604 19628 30660
rect 19684 30604 26908 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 13458 30492 13468 30548
rect 13524 30492 14028 30548
rect 14084 30492 14094 30548
rect 16146 30492 16156 30548
rect 16212 30492 21644 30548
rect 21700 30492 22652 30548
rect 22708 30492 22718 30548
rect 34150 30492 34188 30548
rect 34244 30492 34254 30548
rect 6514 30380 6524 30436
rect 6580 30380 13244 30436
rect 13300 30380 13580 30436
rect 13636 30380 13646 30436
rect 14242 30380 14252 30436
rect 14308 30380 15036 30436
rect 15092 30380 16044 30436
rect 16100 30380 16110 30436
rect 19506 30380 19516 30436
rect 19572 30380 20524 30436
rect 20580 30380 24108 30436
rect 24164 30380 24174 30436
rect 24434 30380 24444 30436
rect 24500 30380 25228 30436
rect 25284 30380 25294 30436
rect 28252 30380 33628 30436
rect 33684 30380 34748 30436
rect 34804 30380 37548 30436
rect 37604 30380 37614 30436
rect 0 30324 800 30352
rect 28252 30324 28308 30380
rect 49200 30324 50000 30352
rect 0 30268 1932 30324
rect 1988 30268 1998 30324
rect 7970 30268 7980 30324
rect 8036 30268 8316 30324
rect 8372 30268 8764 30324
rect 8820 30268 8830 30324
rect 9202 30268 9212 30324
rect 9268 30268 9772 30324
rect 9828 30268 9838 30324
rect 10210 30268 10220 30324
rect 10276 30268 13916 30324
rect 13972 30268 13982 30324
rect 19170 30268 19180 30324
rect 19236 30268 19740 30324
rect 19796 30268 19806 30324
rect 20402 30268 20412 30324
rect 20468 30268 28308 30324
rect 28466 30268 28476 30324
rect 28532 30268 31836 30324
rect 31892 30268 31902 30324
rect 35522 30268 35532 30324
rect 35588 30268 42028 30324
rect 42084 30268 42094 30324
rect 48178 30268 48188 30324
rect 48244 30268 50000 30324
rect 0 30240 800 30268
rect 49200 30240 50000 30268
rect 10322 30156 10332 30212
rect 10388 30156 11788 30212
rect 11844 30156 11854 30212
rect 13010 30156 13020 30212
rect 13076 30156 14252 30212
rect 14308 30156 14700 30212
rect 14756 30156 15036 30212
rect 15092 30156 15932 30212
rect 15988 30156 15998 30212
rect 16706 30156 16716 30212
rect 16772 30156 18060 30212
rect 18116 30156 18126 30212
rect 24546 30156 24556 30212
rect 24612 30156 26012 30212
rect 26068 30156 27692 30212
rect 27748 30156 27758 30212
rect 31154 30156 31164 30212
rect 31220 30156 33068 30212
rect 33124 30156 34412 30212
rect 34468 30156 34478 30212
rect 34636 30156 37212 30212
rect 37268 30156 37278 30212
rect 34636 30100 34692 30156
rect 11330 30044 11340 30100
rect 11396 30044 13132 30100
rect 13188 30044 13198 30100
rect 15138 30044 15148 30100
rect 15204 30044 15708 30100
rect 15764 30044 15774 30100
rect 18946 30044 18956 30100
rect 19012 30044 20188 30100
rect 20244 30044 20636 30100
rect 20692 30044 20702 30100
rect 30706 30044 30716 30100
rect 30772 30044 34692 30100
rect 35746 30044 35756 30100
rect 35812 30044 39676 30100
rect 39732 30044 39742 30100
rect 8866 29932 8876 29988
rect 8932 29932 14476 29988
rect 14532 29932 14542 29988
rect 17826 29932 17836 29988
rect 17892 29932 19180 29988
rect 19236 29932 19246 29988
rect 19628 29932 20076 29988
rect 20132 29932 24668 29988
rect 24724 29932 24734 29988
rect 37090 29932 37100 29988
rect 37156 29932 38556 29988
rect 38612 29932 38892 29988
rect 38948 29932 38958 29988
rect 19628 29876 19684 29932
rect 1474 29820 1484 29876
rect 1540 29820 14812 29876
rect 14868 29820 14878 29876
rect 18946 29820 18956 29876
rect 19012 29820 19684 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 16370 29708 16380 29764
rect 16436 29708 18508 29764
rect 18564 29708 19404 29764
rect 19460 29708 19470 29764
rect 10220 29596 15148 29652
rect 16034 29596 16044 29652
rect 16100 29596 16716 29652
rect 16772 29596 16782 29652
rect 17378 29596 17388 29652
rect 17444 29596 27524 29652
rect 27682 29596 27692 29652
rect 27748 29596 28476 29652
rect 28532 29596 30940 29652
rect 30996 29596 31006 29652
rect 10220 29540 10276 29596
rect 15092 29540 15148 29596
rect 27468 29540 27524 29596
rect 10210 29484 10220 29540
rect 10276 29484 10286 29540
rect 11778 29484 11788 29540
rect 11844 29484 12348 29540
rect 12404 29484 13692 29540
rect 13748 29484 13758 29540
rect 15092 29484 27412 29540
rect 27468 29484 31276 29540
rect 31332 29484 31342 29540
rect 34626 29484 34636 29540
rect 34692 29484 35420 29540
rect 35476 29484 35486 29540
rect 15810 29372 15820 29428
rect 15876 29372 19628 29428
rect 19684 29372 19694 29428
rect 27356 29316 27412 29484
rect 16482 29260 16492 29316
rect 16548 29260 17612 29316
rect 17668 29260 17948 29316
rect 18004 29260 18956 29316
rect 19012 29260 19022 29316
rect 19506 29260 19516 29316
rect 19572 29260 20412 29316
rect 20468 29260 21084 29316
rect 21140 29260 21150 29316
rect 26674 29260 26684 29316
rect 26740 29260 26908 29316
rect 27356 29260 35980 29316
rect 36036 29260 36046 29316
rect 26852 29204 26908 29260
rect 19366 29148 19404 29204
rect 19460 29148 19470 29204
rect 19618 29148 19628 29204
rect 19684 29148 19722 29204
rect 26852 29148 33180 29204
rect 33236 29148 33246 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 18722 28924 18732 28980
rect 18788 28924 19292 28980
rect 19348 28924 19358 28980
rect 4162 28812 4172 28868
rect 4228 28812 8988 28868
rect 9044 28812 9054 28868
rect 9538 28812 9548 28868
rect 9604 28812 18172 28868
rect 18228 28812 18238 28868
rect 0 28756 800 28784
rect 0 28700 1932 28756
rect 1988 28700 1998 28756
rect 2146 28700 2156 28756
rect 2212 28700 4284 28756
rect 4340 28700 7532 28756
rect 7588 28700 7598 28756
rect 16258 28700 16268 28756
rect 16324 28700 38780 28756
rect 38836 28700 39564 28756
rect 39620 28700 39630 28756
rect 0 28672 800 28700
rect 7634 28588 7644 28644
rect 7700 28588 9100 28644
rect 9156 28588 9166 28644
rect 9314 28588 9324 28644
rect 9380 28588 9996 28644
rect 10052 28588 10062 28644
rect 15474 28588 15484 28644
rect 15540 28588 16380 28644
rect 16436 28588 16446 28644
rect 18050 28588 18060 28644
rect 18116 28588 18956 28644
rect 19012 28588 19022 28644
rect 26450 28588 26460 28644
rect 26516 28588 26908 28644
rect 26964 28588 27244 28644
rect 27300 28588 27310 28644
rect 27906 28588 27916 28644
rect 27972 28588 29708 28644
rect 29764 28588 34860 28644
rect 34916 28588 34926 28644
rect 8754 28476 8764 28532
rect 8820 28476 8988 28532
rect 9044 28476 9054 28532
rect 11330 28476 11340 28532
rect 11396 28476 26908 28532
rect 32162 28476 32172 28532
rect 32228 28476 34748 28532
rect 34804 28476 34814 28532
rect 26852 28420 26908 28476
rect 13122 28364 13132 28420
rect 13188 28364 14028 28420
rect 14084 28364 14094 28420
rect 15026 28364 15036 28420
rect 15092 28364 15932 28420
rect 15988 28364 15998 28420
rect 16594 28364 16604 28420
rect 16660 28364 17388 28420
rect 17444 28364 17454 28420
rect 18498 28364 18508 28420
rect 18564 28364 19292 28420
rect 19348 28364 19358 28420
rect 19628 28364 21756 28420
rect 21812 28364 22316 28420
rect 22372 28364 22382 28420
rect 26226 28364 26236 28420
rect 26292 28364 26684 28420
rect 26740 28364 26750 28420
rect 26852 28364 31948 28420
rect 32004 28364 32396 28420
rect 32452 28364 32462 28420
rect 13682 28252 13692 28308
rect 13748 28252 17836 28308
rect 17892 28252 18844 28308
rect 18900 28252 18910 28308
rect 19628 28196 19684 28364
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 17042 28140 17052 28196
rect 17108 28140 17388 28196
rect 17444 28140 17454 28196
rect 17612 28140 19684 28196
rect 17612 28084 17668 28140
rect 5058 28028 5068 28084
rect 5124 28028 9436 28084
rect 9492 28028 9502 28084
rect 9772 28028 17668 28084
rect 18498 28028 18508 28084
rect 18564 28028 33628 28084
rect 33684 28028 33694 28084
rect 8082 27916 8092 27972
rect 8148 27916 9548 27972
rect 9604 27916 9614 27972
rect 9772 27860 9828 28028
rect 16370 27916 16380 27972
rect 16436 27916 16828 27972
rect 16884 27916 17948 27972
rect 18004 27916 18284 27972
rect 18340 27916 18350 27972
rect 19842 27916 19852 27972
rect 19908 27916 20412 27972
rect 20468 27916 34412 27972
rect 34468 27916 34478 27972
rect 3332 27804 4060 27860
rect 4116 27804 7644 27860
rect 7700 27804 7710 27860
rect 8530 27804 8540 27860
rect 8596 27804 8876 27860
rect 8932 27804 8942 27860
rect 9426 27804 9436 27860
rect 9492 27804 9828 27860
rect 14802 27804 14812 27860
rect 14868 27804 14878 27860
rect 17490 27804 17500 27860
rect 17556 27804 20524 27860
rect 20580 27804 20590 27860
rect 20748 27804 27580 27860
rect 27636 27804 30268 27860
rect 30324 27804 30334 27860
rect 40226 27804 40236 27860
rect 40292 27804 41916 27860
rect 41972 27804 41982 27860
rect 3332 27636 3388 27804
rect 14812 27748 14868 27804
rect 20748 27748 20804 27804
rect 7746 27692 7756 27748
rect 7812 27692 9772 27748
rect 9828 27692 9838 27748
rect 14812 27692 16716 27748
rect 16772 27692 16782 27748
rect 19954 27692 19964 27748
rect 20020 27692 20804 27748
rect 20972 27692 29372 27748
rect 29428 27692 29932 27748
rect 29988 27692 31836 27748
rect 31892 27692 31902 27748
rect 32498 27692 32508 27748
rect 32564 27692 33852 27748
rect 33908 27692 33918 27748
rect 34962 27692 34972 27748
rect 35028 27692 35980 27748
rect 36036 27692 36046 27748
rect 2930 27580 2940 27636
rect 2996 27580 3388 27636
rect 4274 27580 4284 27636
rect 4340 27580 8204 27636
rect 8260 27580 8270 27636
rect 8530 27580 8540 27636
rect 8596 27580 9884 27636
rect 9940 27580 9950 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 20972 27412 21028 27692
rect 23426 27580 23436 27636
rect 23492 27580 23996 27636
rect 24052 27580 24062 27636
rect 21298 27468 21308 27524
rect 21364 27468 30156 27524
rect 30212 27468 30222 27524
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 11554 27356 11564 27412
rect 11620 27356 21028 27412
rect 24098 27356 24108 27412
rect 24164 27356 34356 27412
rect 6850 27244 6860 27300
rect 6916 27244 8316 27300
rect 8372 27244 8382 27300
rect 15810 27244 15820 27300
rect 15876 27244 17500 27300
rect 17556 27244 18396 27300
rect 18452 27244 18462 27300
rect 19394 27244 19404 27300
rect 19460 27244 19964 27300
rect 20020 27244 20030 27300
rect 20514 27244 20524 27300
rect 20580 27244 21308 27300
rect 21364 27244 21374 27300
rect 22306 27244 22316 27300
rect 22372 27244 23100 27300
rect 23156 27244 23166 27300
rect 26226 27244 26236 27300
rect 26292 27244 26908 27300
rect 26964 27244 27356 27300
rect 27412 27244 27422 27300
rect 0 27188 800 27216
rect 0 27132 1932 27188
rect 1988 27132 1998 27188
rect 16594 27132 16604 27188
rect 16660 27132 19292 27188
rect 19348 27132 19358 27188
rect 22316 27132 23436 27188
rect 23492 27132 23884 27188
rect 23940 27132 23950 27188
rect 26338 27132 26348 27188
rect 26404 27132 27468 27188
rect 27524 27132 27534 27188
rect 31938 27132 31948 27188
rect 32004 27132 32396 27188
rect 32452 27132 32462 27188
rect 0 27104 800 27132
rect 22316 27076 22372 27132
rect 34300 27076 34356 27356
rect 9986 27020 9996 27076
rect 10052 27020 10444 27076
rect 10500 27020 10510 27076
rect 18162 27020 18172 27076
rect 18228 27020 20412 27076
rect 20468 27020 21196 27076
rect 21252 27020 21262 27076
rect 21634 27020 21644 27076
rect 21700 27020 21980 27076
rect 22036 27020 22046 27076
rect 22306 27020 22316 27076
rect 22372 27020 22382 27076
rect 23314 27020 23324 27076
rect 23380 27020 24108 27076
rect 24164 27020 24174 27076
rect 25218 27020 25228 27076
rect 25284 27020 25900 27076
rect 25956 27020 25966 27076
rect 34300 27020 35532 27076
rect 35588 27020 36316 27076
rect 36372 27020 36382 27076
rect 36316 26964 36372 27020
rect 2146 26908 2156 26964
rect 2212 26908 4508 26964
rect 4564 26908 6748 26964
rect 6804 26908 6814 26964
rect 18610 26908 18620 26964
rect 18676 26908 19292 26964
rect 19348 26908 19358 26964
rect 23874 26908 23884 26964
rect 23940 26908 24892 26964
rect 24948 26908 25676 26964
rect 25732 26908 25742 26964
rect 36316 26908 40236 26964
rect 40292 26908 40302 26964
rect 7410 26796 7420 26852
rect 7476 26796 9100 26852
rect 9156 26796 9166 26852
rect 10210 26796 10220 26852
rect 10276 26796 14364 26852
rect 14420 26796 14430 26852
rect 15092 26796 16940 26852
rect 16996 26796 17006 26852
rect 19170 26796 19180 26852
rect 19236 26796 20300 26852
rect 20356 26796 20366 26852
rect 21970 26796 21980 26852
rect 22036 26796 22988 26852
rect 23044 26796 23054 26852
rect 23762 26796 23772 26852
rect 23828 26796 24108 26852
rect 24164 26796 24174 26852
rect 25330 26796 25340 26852
rect 25396 26796 26572 26852
rect 26628 26796 26638 26852
rect 33506 26796 33516 26852
rect 33572 26796 36204 26852
rect 36260 26796 37100 26852
rect 37156 26796 38556 26852
rect 38612 26796 38622 26852
rect 15092 26740 15148 26796
rect 8754 26684 8764 26740
rect 8820 26684 15148 26740
rect 16370 26684 16380 26740
rect 16436 26684 17612 26740
rect 17668 26684 18508 26740
rect 18564 26684 18574 26740
rect 34514 26684 34524 26740
rect 34580 26684 35868 26740
rect 35924 26684 35934 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 21746 26572 21756 26628
rect 21812 26572 22876 26628
rect 22932 26572 22942 26628
rect 1586 26460 1596 26516
rect 1652 26460 3388 26516
rect 13010 26460 13020 26516
rect 13076 26460 14700 26516
rect 14756 26460 14766 26516
rect 16706 26460 16716 26516
rect 16772 26460 19964 26516
rect 20020 26460 20030 26516
rect 20290 26460 20300 26516
rect 20356 26460 21532 26516
rect 21588 26460 21598 26516
rect 22530 26460 22540 26516
rect 22596 26460 24332 26516
rect 24388 26460 25004 26516
rect 25060 26460 25070 26516
rect 34402 26460 34412 26516
rect 34468 26460 36428 26516
rect 36484 26460 36494 26516
rect 3332 26404 3388 26460
rect 3332 26348 16044 26404
rect 16100 26348 16268 26404
rect 16324 26348 16334 26404
rect 18956 26348 25452 26404
rect 25508 26348 26796 26404
rect 26852 26348 26862 26404
rect 18956 26292 19012 26348
rect 14018 26236 14028 26292
rect 14084 26236 14588 26292
rect 14644 26236 15260 26292
rect 15316 26236 15326 26292
rect 18946 26236 18956 26292
rect 19012 26236 19022 26292
rect 19842 26236 19852 26292
rect 19908 26236 19918 26292
rect 21410 26236 21420 26292
rect 21476 26236 21980 26292
rect 22036 26236 29484 26292
rect 29540 26236 31612 26292
rect 31668 26236 31678 26292
rect 4946 26124 4956 26180
rect 5012 26124 8092 26180
rect 8148 26124 8158 26180
rect 17266 26124 17276 26180
rect 17332 26124 18172 26180
rect 18228 26124 18238 26180
rect 19852 26068 19908 26236
rect 20178 26124 20188 26180
rect 20244 26124 21196 26180
rect 21252 26124 33404 26180
rect 33460 26124 33470 26180
rect 36866 26124 36876 26180
rect 36932 26124 37996 26180
rect 38052 26124 38062 26180
rect 8418 26012 8428 26068
rect 8484 26012 9212 26068
rect 9268 26012 9278 26068
rect 9958 26012 9996 26068
rect 10052 26012 10062 26068
rect 10658 26012 10668 26068
rect 10724 26012 19908 26068
rect 22082 26012 22092 26068
rect 22148 26012 22876 26068
rect 22932 26012 23100 26068
rect 23156 26012 23166 26068
rect 23426 26012 23436 26068
rect 23492 26012 24108 26068
rect 24164 26012 24174 26068
rect 38612 26012 39340 26068
rect 39396 26012 39406 26068
rect 23100 25956 23156 26012
rect 14690 25900 14700 25956
rect 14756 25900 16996 25956
rect 17714 25900 17724 25956
rect 17780 25900 21868 25956
rect 21924 25900 21934 25956
rect 23100 25900 25340 25956
rect 25396 25900 25406 25956
rect 33506 25900 33516 25956
rect 33572 25900 34636 25956
rect 34692 25900 34702 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 7410 25788 7420 25844
rect 7476 25788 7980 25844
rect 8036 25788 8046 25844
rect 15810 25788 15820 25844
rect 15876 25788 16716 25844
rect 16772 25788 16782 25844
rect 16940 25732 16996 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 23650 25788 23660 25844
rect 23716 25788 25228 25844
rect 25284 25788 25294 25844
rect 30716 25788 32844 25844
rect 32900 25788 33628 25844
rect 33684 25788 34300 25844
rect 34356 25788 34366 25844
rect 30716 25732 30772 25788
rect 38612 25732 38668 26012
rect 6850 25676 6860 25732
rect 6916 25676 8204 25732
rect 8260 25676 8270 25732
rect 15922 25676 15932 25732
rect 15988 25676 16604 25732
rect 16660 25676 16670 25732
rect 16902 25676 16940 25732
rect 16996 25676 17612 25732
rect 17668 25676 17678 25732
rect 23426 25676 23436 25732
rect 23492 25676 30772 25732
rect 30828 25676 38668 25732
rect 0 25620 800 25648
rect 30828 25620 30884 25676
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 12002 25564 12012 25620
rect 12068 25564 14924 25620
rect 14980 25564 14990 25620
rect 15708 25564 16492 25620
rect 16548 25564 30884 25620
rect 32386 25564 32396 25620
rect 32452 25564 33292 25620
rect 33348 25564 33358 25620
rect 34748 25564 35084 25620
rect 35140 25564 35756 25620
rect 35812 25564 40012 25620
rect 40068 25564 40078 25620
rect 0 25536 800 25564
rect 15708 25396 15764 25564
rect 34748 25508 34804 25564
rect 20738 25452 20748 25508
rect 20804 25452 22372 25508
rect 22316 25396 22372 25452
rect 26852 25452 34804 25508
rect 34962 25452 34972 25508
rect 35028 25452 38892 25508
rect 38948 25452 38958 25508
rect 39330 25452 39340 25508
rect 39396 25452 40124 25508
rect 40180 25452 40190 25508
rect 42018 25452 42028 25508
rect 42084 25452 47852 25508
rect 47908 25452 47918 25508
rect 26852 25396 26908 25452
rect 40124 25396 40180 25452
rect 13906 25340 13916 25396
rect 13972 25340 14252 25396
rect 14308 25340 14812 25396
rect 14868 25340 14878 25396
rect 15026 25340 15036 25396
rect 15092 25340 15764 25396
rect 15922 25340 15932 25396
rect 15988 25340 18620 25396
rect 18676 25340 18686 25396
rect 22306 25340 22316 25396
rect 22372 25340 26908 25396
rect 33394 25340 33404 25396
rect 33460 25340 34188 25396
rect 34244 25340 34524 25396
rect 34580 25340 34590 25396
rect 34850 25340 34860 25396
rect 34916 25340 36316 25396
rect 36372 25340 36382 25396
rect 40124 25340 43372 25396
rect 43428 25340 43438 25396
rect 8642 25228 8652 25284
rect 8708 25228 18396 25284
rect 18452 25228 18462 25284
rect 19628 25228 19740 25284
rect 19796 25228 19806 25284
rect 26786 25228 26796 25284
rect 26852 25228 27244 25284
rect 27300 25228 45052 25284
rect 45108 25228 45118 25284
rect 47618 25228 47628 25284
rect 47684 25228 48188 25284
rect 48244 25228 48254 25284
rect 19628 25172 19684 25228
rect 7746 25116 7756 25172
rect 7812 25116 8316 25172
rect 8372 25116 8382 25172
rect 15250 25116 15260 25172
rect 15316 25116 15484 25172
rect 15540 25116 15550 25172
rect 18498 25116 18508 25172
rect 18564 25116 19684 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 14242 25004 14252 25060
rect 14308 25004 14924 25060
rect 14980 25004 14990 25060
rect 16482 25004 16492 25060
rect 16548 25004 17164 25060
rect 17220 25004 17230 25060
rect 19058 25004 19068 25060
rect 19124 25004 19292 25060
rect 19348 25004 19358 25060
rect 34262 25004 34300 25060
rect 34356 25004 34366 25060
rect 49200 24948 50000 24976
rect 6402 24892 6412 24948
rect 6468 24892 17612 24948
rect 17668 24892 17948 24948
rect 18004 24892 18014 24948
rect 20402 24892 20412 24948
rect 20468 24892 20860 24948
rect 20916 24892 20926 24948
rect 34402 24892 34412 24948
rect 34468 24892 34478 24948
rect 48178 24892 48188 24948
rect 48244 24892 50000 24948
rect 34412 24836 34468 24892
rect 49200 24864 50000 24892
rect 8166 24780 8204 24836
rect 8260 24780 8270 24836
rect 8978 24780 8988 24836
rect 9044 24780 13916 24836
rect 13972 24780 13982 24836
rect 15474 24780 15484 24836
rect 15540 24780 18844 24836
rect 18900 24780 19852 24836
rect 19908 24780 19918 24836
rect 22866 24780 22876 24836
rect 22932 24780 23996 24836
rect 24052 24780 26348 24836
rect 26404 24780 26414 24836
rect 26786 24780 26796 24836
rect 26852 24780 30324 24836
rect 33842 24780 33852 24836
rect 33908 24780 34748 24836
rect 34804 24780 34814 24836
rect 11106 24668 11116 24724
rect 11172 24668 11788 24724
rect 11844 24668 12236 24724
rect 12292 24668 12796 24724
rect 12852 24668 12862 24724
rect 16706 24668 16716 24724
rect 16772 24668 18620 24724
rect 18676 24668 18686 24724
rect 30268 24612 30324 24780
rect 30482 24668 30492 24724
rect 30548 24668 31052 24724
rect 31108 24668 36428 24724
rect 36484 24668 36494 24724
rect 36866 24668 36876 24724
rect 36932 24668 39676 24724
rect 39732 24668 39742 24724
rect 2818 24556 2828 24612
rect 2884 24556 4284 24612
rect 4340 24556 4350 24612
rect 9874 24556 9884 24612
rect 9940 24556 14812 24612
rect 14868 24556 16156 24612
rect 16212 24556 16222 24612
rect 16370 24556 16380 24612
rect 16436 24556 18284 24612
rect 18340 24556 18350 24612
rect 18498 24556 18508 24612
rect 18564 24556 19180 24612
rect 19236 24556 19246 24612
rect 30268 24556 34076 24612
rect 34132 24556 34860 24612
rect 34916 24556 34926 24612
rect 8866 24444 8876 24500
rect 8932 24444 11676 24500
rect 11732 24444 11742 24500
rect 16594 24444 16604 24500
rect 16660 24444 17276 24500
rect 17332 24444 17342 24500
rect 33590 24444 33628 24500
rect 33684 24444 33694 24500
rect 36642 24444 36652 24500
rect 36708 24444 37772 24500
rect 37828 24444 37838 24500
rect 39778 24444 39788 24500
rect 39844 24444 41244 24500
rect 41300 24444 41310 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 23986 24220 23996 24276
rect 24052 24220 24556 24276
rect 24612 24220 24622 24276
rect 34374 24220 34412 24276
rect 34468 24220 34478 24276
rect 12450 24108 12460 24164
rect 12516 24108 13580 24164
rect 13636 24108 13646 24164
rect 34066 24108 34076 24164
rect 34132 24108 34300 24164
rect 34356 24108 34366 24164
rect 0 24052 800 24080
rect 0 23996 1932 24052
rect 1988 23996 1998 24052
rect 7634 23996 7644 24052
rect 7700 23996 8764 24052
rect 8820 23996 9772 24052
rect 9828 23996 28588 24052
rect 28644 23996 29148 24052
rect 29204 23996 30828 24052
rect 30884 23996 30894 24052
rect 0 23968 800 23996
rect 30828 23940 30884 23996
rect 4274 23884 4284 23940
rect 4340 23884 6748 23940
rect 6804 23884 6814 23940
rect 7858 23884 7868 23940
rect 7924 23884 10668 23940
rect 10724 23884 10734 23940
rect 27570 23884 27580 23940
rect 27636 23884 29484 23940
rect 29540 23884 29550 23940
rect 30828 23884 31500 23940
rect 31556 23884 31566 23940
rect 36418 23884 36428 23940
rect 36484 23884 37100 23940
rect 37156 23884 37884 23940
rect 37940 23884 40124 23940
rect 40180 23884 40460 23940
rect 40516 23884 40526 23940
rect 11666 23772 11676 23828
rect 11732 23772 11900 23828
rect 11956 23772 12684 23828
rect 12740 23772 12750 23828
rect 13570 23772 13580 23828
rect 13636 23772 14028 23828
rect 14084 23772 14094 23828
rect 14578 23772 14588 23828
rect 14644 23772 16492 23828
rect 16548 23772 16558 23828
rect 19170 23772 19180 23828
rect 19236 23772 20188 23828
rect 20244 23772 20254 23828
rect 23314 23772 23324 23828
rect 23380 23772 23772 23828
rect 23828 23772 24668 23828
rect 24724 23772 24734 23828
rect 25554 23772 25564 23828
rect 25620 23772 29596 23828
rect 29652 23772 29662 23828
rect 12684 23716 12740 23772
rect 12684 23660 15148 23716
rect 17154 23660 17164 23716
rect 17220 23660 22764 23716
rect 22820 23660 22830 23716
rect 15092 23604 15148 23660
rect 5954 23548 5964 23604
rect 6020 23548 7420 23604
rect 7476 23548 7486 23604
rect 12674 23548 12684 23604
rect 12740 23548 14588 23604
rect 14644 23548 14654 23604
rect 15092 23548 17388 23604
rect 17444 23548 17454 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 21298 23436 21308 23492
rect 21364 23436 23324 23492
rect 23380 23436 24668 23492
rect 24724 23436 25228 23492
rect 25284 23436 25294 23492
rect 3332 23324 8036 23380
rect 17266 23324 17276 23380
rect 17332 23324 17948 23380
rect 18004 23324 18014 23380
rect 18162 23324 18172 23380
rect 18228 23324 18844 23380
rect 18900 23324 18910 23380
rect 20850 23324 20860 23380
rect 20916 23324 28308 23380
rect 3332 23268 3388 23324
rect 3154 23212 3164 23268
rect 3220 23212 3388 23268
rect 4274 23212 4284 23268
rect 4340 23212 5740 23268
rect 5796 23212 5806 23268
rect 4284 23156 4340 23212
rect 7980 23156 8036 23324
rect 13570 23212 13580 23268
rect 13636 23212 13646 23268
rect 15092 23212 15260 23268
rect 15316 23212 15326 23268
rect 16146 23212 16156 23268
rect 16212 23212 21532 23268
rect 21588 23212 21598 23268
rect 21858 23212 21868 23268
rect 21924 23212 22204 23268
rect 22260 23212 26908 23268
rect 13580 23156 13636 23212
rect 15092 23156 15148 23212
rect 2034 23100 2044 23156
rect 2100 23100 4340 23156
rect 5842 23100 5852 23156
rect 5908 23100 7308 23156
rect 7364 23100 7374 23156
rect 7970 23100 7980 23156
rect 8036 23100 8046 23156
rect 13580 23100 15148 23156
rect 16370 23100 16380 23156
rect 16436 23100 17500 23156
rect 17556 23100 17566 23156
rect 17714 23100 17724 23156
rect 17780 23100 17948 23156
rect 18004 23100 18014 23156
rect 26852 23044 26908 23212
rect 28252 23156 28308 23324
rect 27682 23100 27692 23156
rect 27748 23100 28028 23156
rect 28084 23100 28094 23156
rect 28242 23100 28252 23156
rect 28308 23100 30828 23156
rect 30884 23100 30894 23156
rect 5170 22988 5180 23044
rect 5236 22988 6300 23044
rect 6356 22988 6366 23044
rect 7746 22988 7756 23044
rect 7812 22988 8316 23044
rect 8372 22988 8382 23044
rect 12226 22988 12236 23044
rect 12292 22988 14028 23044
rect 14084 22988 14094 23044
rect 20290 22988 20300 23044
rect 20356 22988 21084 23044
rect 21140 22988 21150 23044
rect 26852 22988 28812 23044
rect 28868 22988 29708 23044
rect 29764 22988 30268 23044
rect 30324 22988 33180 23044
rect 33236 22988 33246 23044
rect 7074 22764 7084 22820
rect 7140 22764 9436 22820
rect 9492 22764 9502 22820
rect 15250 22764 15260 22820
rect 15316 22764 15820 22820
rect 15876 22764 15886 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 9090 22652 9100 22708
rect 9156 22652 22428 22708
rect 22484 22652 23772 22708
rect 23828 22652 23838 22708
rect 4498 22540 4508 22596
rect 4564 22540 7644 22596
rect 7700 22540 7710 22596
rect 15092 22540 15708 22596
rect 15764 22540 15774 22596
rect 0 22484 800 22512
rect 15092 22484 15148 22540
rect 0 22428 1932 22484
rect 1988 22428 1998 22484
rect 4162 22428 4172 22484
rect 4228 22428 7196 22484
rect 7252 22428 7262 22484
rect 14354 22428 14364 22484
rect 14420 22428 15148 22484
rect 15558 22428 15596 22484
rect 15652 22428 15662 22484
rect 18722 22428 18732 22484
rect 18788 22428 19404 22484
rect 19460 22428 19470 22484
rect 0 22400 800 22428
rect 14018 22316 14028 22372
rect 14084 22316 15148 22372
rect 15092 22260 15148 22316
rect 6626 22204 6636 22260
rect 6692 22204 8764 22260
rect 8820 22204 8830 22260
rect 9986 22204 9996 22260
rect 10052 22204 13580 22260
rect 13636 22204 13646 22260
rect 15092 22204 17948 22260
rect 18004 22204 18014 22260
rect 7522 22092 7532 22148
rect 7588 22092 8316 22148
rect 8372 22092 8382 22148
rect 12002 22092 12012 22148
rect 12068 22092 13804 22148
rect 13860 22092 14700 22148
rect 14756 22092 15148 22148
rect 16706 22092 16716 22148
rect 16772 22092 18060 22148
rect 18116 22092 18284 22148
rect 18340 22092 18350 22148
rect 20850 22092 20860 22148
rect 20916 22092 21308 22148
rect 21364 22092 22204 22148
rect 22260 22092 22270 22148
rect 23090 22092 23100 22148
rect 23156 22092 23660 22148
rect 23716 22092 24668 22148
rect 24724 22092 24734 22148
rect 25554 22092 25564 22148
rect 25620 22092 27468 22148
rect 27524 22092 29596 22148
rect 29652 22092 30044 22148
rect 30100 22092 34188 22148
rect 34244 22092 34254 22148
rect 15092 22036 15148 22092
rect 10098 21980 10108 22036
rect 10164 21980 10174 22036
rect 15092 21980 15372 22036
rect 15428 21980 15438 22036
rect 10108 21812 10164 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 11890 21868 11900 21924
rect 11956 21868 16044 21924
rect 16100 21868 16110 21924
rect 20738 21868 20748 21924
rect 20804 21868 21756 21924
rect 21812 21868 21822 21924
rect 25218 21868 25228 21924
rect 25284 21868 25294 21924
rect 26114 21868 26124 21924
rect 26180 21868 30044 21924
rect 30100 21868 30110 21924
rect 25228 21812 25284 21868
rect 10108 21756 11452 21812
rect 11508 21756 11518 21812
rect 12226 21756 12236 21812
rect 12292 21756 13468 21812
rect 13524 21756 15148 21812
rect 15204 21756 15708 21812
rect 15764 21756 15774 21812
rect 16706 21756 16716 21812
rect 16772 21756 19068 21812
rect 19124 21756 22204 21812
rect 22260 21756 24668 21812
rect 24724 21756 25284 21812
rect 31714 21756 31724 21812
rect 31780 21756 34412 21812
rect 34468 21756 35196 21812
rect 35252 21756 38668 21812
rect 8978 21644 8988 21700
rect 9044 21644 11564 21700
rect 11620 21644 11630 21700
rect 19842 21644 19852 21700
rect 19908 21644 20748 21700
rect 20804 21644 20814 21700
rect 21644 21644 22876 21700
rect 22932 21644 22942 21700
rect 25330 21644 25340 21700
rect 25396 21644 25900 21700
rect 25956 21644 25966 21700
rect 21644 21588 21700 21644
rect 38612 21588 38668 21756
rect 9650 21532 9660 21588
rect 9716 21532 10108 21588
rect 10164 21532 10174 21588
rect 10658 21532 10668 21588
rect 10724 21532 12124 21588
rect 12180 21532 12190 21588
rect 14466 21532 14476 21588
rect 14532 21532 19404 21588
rect 19460 21532 19470 21588
rect 21634 21532 21644 21588
rect 21700 21532 21710 21588
rect 22530 21532 22540 21588
rect 22596 21532 22988 21588
rect 23044 21532 23212 21588
rect 23268 21532 23660 21588
rect 23716 21532 23726 21588
rect 24322 21532 24332 21588
rect 24388 21532 25116 21588
rect 25172 21532 32060 21588
rect 32116 21532 34748 21588
rect 34804 21532 35420 21588
rect 35476 21532 35486 21588
rect 38612 21532 46284 21588
rect 46340 21532 46350 21588
rect 7634 21420 7644 21476
rect 7700 21420 8428 21476
rect 8484 21420 8494 21476
rect 15586 21420 15596 21476
rect 15652 21420 18396 21476
rect 18452 21420 18462 21476
rect 20514 21420 20524 21476
rect 20580 21420 21084 21476
rect 21140 21420 21150 21476
rect 24770 21420 24780 21476
rect 24836 21420 25340 21476
rect 25396 21420 25406 21476
rect 16370 21308 16380 21364
rect 16436 21308 23436 21364
rect 23492 21308 23502 21364
rect 8978 21196 8988 21252
rect 9044 21196 12572 21252
rect 12628 21196 14924 21252
rect 14980 21196 14990 21252
rect 16146 21196 16156 21252
rect 16212 21196 16604 21252
rect 16660 21196 16670 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 14102 21084 14140 21140
rect 14196 21084 14206 21140
rect 12898 20972 12908 21028
rect 12964 20972 14588 21028
rect 14644 20972 14654 21028
rect 0 20916 800 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 10882 20860 10892 20916
rect 10948 20860 12348 20916
rect 12404 20860 12796 20916
rect 12852 20860 15596 20916
rect 15652 20860 15662 20916
rect 23874 20860 23884 20916
rect 23940 20860 24220 20916
rect 24276 20860 24556 20916
rect 24612 20860 25564 20916
rect 25620 20860 25630 20916
rect 33842 20860 33852 20916
rect 33908 20860 34972 20916
rect 35028 20860 37212 20916
rect 37268 20860 37884 20916
rect 37940 20860 37950 20916
rect 0 20832 800 20860
rect 2258 20748 2268 20804
rect 2324 20748 4284 20804
rect 4340 20748 5852 20804
rect 5908 20748 5918 20804
rect 14354 20748 14364 20804
rect 14420 20748 16268 20804
rect 16324 20748 16334 20804
rect 22530 20748 22540 20804
rect 22596 20748 23324 20804
rect 23380 20748 23390 20804
rect 24994 20748 25004 20804
rect 25060 20748 26236 20804
rect 26292 20748 26302 20804
rect 29362 20748 29372 20804
rect 29428 20748 29932 20804
rect 29988 20748 29998 20804
rect 22540 20692 22596 20748
rect 19954 20636 19964 20692
rect 20020 20636 20412 20692
rect 20468 20636 22596 20692
rect 30146 20636 30156 20692
rect 30212 20636 33068 20692
rect 33124 20636 33134 20692
rect 37426 20636 37436 20692
rect 37492 20636 39004 20692
rect 39060 20636 39070 20692
rect 8306 20524 8316 20580
rect 8372 20524 9100 20580
rect 9156 20524 9436 20580
rect 9492 20524 10052 20580
rect 9996 20468 10052 20524
rect 14364 20524 17276 20580
rect 17332 20524 25004 20580
rect 25060 20524 25070 20580
rect 35746 20524 35756 20580
rect 35812 20524 36652 20580
rect 36708 20524 36718 20580
rect 14364 20468 14420 20524
rect 9986 20412 9996 20468
rect 10052 20412 10062 20468
rect 14354 20412 14364 20468
rect 14420 20412 14430 20468
rect 14578 20412 14588 20468
rect 14644 20412 15148 20468
rect 15204 20412 16156 20468
rect 16212 20412 16222 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 21074 20300 21084 20356
rect 21140 20300 21980 20356
rect 22036 20300 22316 20356
rect 22372 20300 37884 20356
rect 37940 20300 37950 20356
rect 15922 20188 15932 20244
rect 15988 20188 16716 20244
rect 16772 20188 16782 20244
rect 30818 20188 30828 20244
rect 30884 20188 31836 20244
rect 31892 20188 31902 20244
rect 35746 20188 35756 20244
rect 35812 20188 37212 20244
rect 37268 20188 37278 20244
rect 39106 20188 39116 20244
rect 39172 20188 39676 20244
rect 39732 20188 39742 20244
rect 13794 20076 13804 20132
rect 13860 20076 15372 20132
rect 15428 20076 15438 20132
rect 15586 20076 15596 20132
rect 15652 20076 24668 20132
rect 24724 20076 25452 20132
rect 25508 20076 25518 20132
rect 26450 20076 26460 20132
rect 26516 20076 27020 20132
rect 27076 20076 27086 20132
rect 30258 20076 30268 20132
rect 30324 20076 30716 20132
rect 30772 20076 30782 20132
rect 33404 20076 35084 20132
rect 35140 20076 35532 20132
rect 35588 20076 35598 20132
rect 46162 20076 46172 20132
rect 46228 20076 47852 20132
rect 47908 20076 47918 20132
rect 33404 20020 33460 20076
rect 10994 19964 11004 20020
rect 11060 19964 11564 20020
rect 11620 19964 11630 20020
rect 18050 19964 18060 20020
rect 18116 19964 21308 20020
rect 21364 19964 22652 20020
rect 22708 19964 22718 20020
rect 23762 19964 23772 20020
rect 23828 19964 26796 20020
rect 26852 19964 33460 20020
rect 35186 19964 35196 20020
rect 35252 19964 36540 20020
rect 36596 19964 36606 20020
rect 1698 19852 1708 19908
rect 1764 19852 2492 19908
rect 2548 19852 2558 19908
rect 7970 19852 7980 19908
rect 8036 19852 8764 19908
rect 8820 19852 8830 19908
rect 10658 19852 10668 19908
rect 10724 19852 11900 19908
rect 11956 19852 12908 19908
rect 12964 19852 12974 19908
rect 25890 19852 25900 19908
rect 25956 19852 31948 19908
rect 32004 19852 34860 19908
rect 34916 19852 35420 19908
rect 35476 19852 35486 19908
rect 36418 19852 36428 19908
rect 36484 19852 37996 19908
rect 38052 19852 38062 19908
rect 39218 19852 39228 19908
rect 39284 19852 40124 19908
rect 40180 19852 40190 19908
rect 2034 19740 2044 19796
rect 2100 19740 15148 19796
rect 24546 19740 24556 19796
rect 24612 19740 30268 19796
rect 30324 19740 30334 19796
rect 30818 19740 30828 19796
rect 30884 19740 31724 19796
rect 31780 19740 31790 19796
rect 15092 19684 15148 19740
rect 8418 19628 8428 19684
rect 8484 19628 9660 19684
rect 9716 19628 9726 19684
rect 12338 19628 12348 19684
rect 12404 19628 13804 19684
rect 13860 19628 13870 19684
rect 15092 19628 20412 19684
rect 20468 19628 20748 19684
rect 20804 19628 22876 19684
rect 22932 19628 22942 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 49200 19572 50000 19600
rect 11330 19516 11340 19572
rect 11396 19516 11900 19572
rect 11956 19516 12796 19572
rect 12852 19516 12862 19572
rect 48178 19516 48188 19572
rect 48244 19516 50000 19572
rect 49200 19488 50000 19516
rect 12562 19404 12572 19460
rect 12628 19404 14028 19460
rect 14084 19404 14094 19460
rect 0 19348 800 19376
rect 0 19292 1708 19348
rect 1764 19292 1774 19348
rect 10658 19292 10668 19348
rect 10724 19292 12348 19348
rect 12404 19292 12414 19348
rect 13010 19292 13020 19348
rect 13076 19292 13804 19348
rect 13860 19292 13870 19348
rect 15250 19292 15260 19348
rect 15316 19292 16380 19348
rect 16436 19292 16446 19348
rect 32162 19292 32172 19348
rect 32228 19292 32844 19348
rect 32900 19292 37212 19348
rect 37268 19292 38108 19348
rect 38164 19292 41132 19348
rect 41188 19292 41198 19348
rect 0 19264 800 19292
rect 3332 19180 8316 19236
rect 8372 19180 8382 19236
rect 9762 19180 9772 19236
rect 9828 19180 12124 19236
rect 12180 19180 13916 19236
rect 13972 19180 13982 19236
rect 29698 19180 29708 19236
rect 29764 19180 30604 19236
rect 30660 19180 30670 19236
rect 34626 19180 34636 19236
rect 34692 19180 35980 19236
rect 36036 19180 36428 19236
rect 36484 19180 36988 19236
rect 37044 19180 37054 19236
rect 3332 19124 3388 19180
rect 1922 19068 1932 19124
rect 1988 19068 3388 19124
rect 7186 19068 7196 19124
rect 7252 19068 21532 19124
rect 21588 19068 25676 19124
rect 25732 19068 26460 19124
rect 26516 19068 26526 19124
rect 2706 18956 2716 19012
rect 2772 18956 8876 19012
rect 8932 18956 11004 19012
rect 11060 18956 11070 19012
rect 27122 18956 27132 19012
rect 27188 18956 27580 19012
rect 27636 18956 27646 19012
rect 30706 18956 30716 19012
rect 30772 18956 31388 19012
rect 31444 18956 33628 19012
rect 33684 18956 33694 19012
rect 35858 18956 35868 19012
rect 35924 18956 36316 19012
rect 36372 18956 39228 19012
rect 39284 18956 39294 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 9650 18620 9660 18676
rect 9716 18620 10724 18676
rect 15138 18620 15148 18676
rect 15204 18620 15596 18676
rect 15652 18620 15662 18676
rect 10668 18564 10724 18620
rect 8866 18508 8876 18564
rect 8932 18508 9772 18564
rect 9828 18508 10108 18564
rect 10164 18508 10174 18564
rect 10658 18508 10668 18564
rect 10724 18508 11564 18564
rect 11620 18508 12012 18564
rect 12068 18508 12078 18564
rect 18162 18508 18172 18564
rect 18228 18508 18620 18564
rect 18676 18508 18686 18564
rect 6514 18396 6524 18452
rect 6580 18396 7196 18452
rect 7252 18396 7262 18452
rect 30482 18396 30492 18452
rect 30548 18396 35868 18452
rect 35924 18396 35934 18452
rect 1698 18284 1708 18340
rect 1764 18284 2492 18340
rect 2548 18284 2558 18340
rect 14802 18284 14812 18340
rect 14868 18284 17612 18340
rect 17668 18284 17948 18340
rect 18004 18284 18014 18340
rect 19394 18284 19404 18340
rect 19460 18284 21420 18340
rect 21476 18284 31388 18340
rect 31444 18284 31836 18340
rect 31892 18284 31902 18340
rect 32722 18284 32732 18340
rect 32788 18284 33292 18340
rect 33348 18284 33358 18340
rect 2034 18172 2044 18228
rect 2100 18172 15148 18228
rect 18050 18172 18060 18228
rect 18116 18172 19516 18228
rect 19572 18172 19582 18228
rect 15092 18116 15148 18172
rect 15092 18060 25340 18116
rect 25396 18060 26124 18116
rect 26180 18060 29036 18116
rect 29092 18060 29820 18116
rect 29876 18060 29886 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 9762 17948 9772 18004
rect 9828 17948 24556 18004
rect 24612 17948 24622 18004
rect 8642 17836 8652 17892
rect 8708 17836 9100 17892
rect 9156 17836 26908 17892
rect 26964 17836 27468 17892
rect 27524 17836 27534 17892
rect 0 17780 800 17808
rect 0 17724 1708 17780
rect 1764 17724 1774 17780
rect 5058 17724 5068 17780
rect 5124 17724 6188 17780
rect 6244 17724 6254 17780
rect 18386 17724 18396 17780
rect 18452 17724 20748 17780
rect 20804 17724 21532 17780
rect 21588 17724 23100 17780
rect 23156 17724 23166 17780
rect 0 17696 800 17724
rect 21298 17612 21308 17668
rect 21364 17612 21644 17668
rect 21700 17612 25676 17668
rect 25732 17612 25742 17668
rect 2930 17500 2940 17556
rect 2996 17500 6748 17556
rect 6804 17500 6814 17556
rect 6962 17500 6972 17556
rect 7028 17500 8428 17556
rect 8484 17500 8494 17556
rect 19058 17500 19068 17556
rect 19124 17500 19740 17556
rect 19796 17500 20300 17556
rect 20356 17500 20366 17556
rect 27570 17500 27580 17556
rect 27636 17500 28140 17556
rect 28196 17500 28206 17556
rect 29362 17500 29372 17556
rect 29428 17500 30380 17556
rect 30436 17500 30716 17556
rect 30772 17500 34412 17556
rect 34468 17500 34478 17556
rect 2258 17388 2268 17444
rect 2324 17388 3388 17444
rect 8194 17388 8204 17444
rect 8260 17388 8540 17444
rect 8596 17388 21980 17444
rect 22036 17388 22046 17444
rect 26002 17388 26012 17444
rect 26068 17388 28588 17444
rect 28644 17388 30604 17444
rect 30660 17388 30670 17444
rect 35858 17388 35868 17444
rect 35924 17388 36092 17444
rect 36148 17388 37100 17444
rect 37156 17388 39116 17444
rect 39172 17388 39900 17444
rect 39956 17388 39966 17444
rect 3332 17220 3388 17388
rect 10994 17276 11004 17332
rect 11060 17276 13804 17332
rect 13860 17276 15708 17332
rect 15764 17276 15774 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 3332 17164 3948 17220
rect 4004 17164 11788 17220
rect 11844 17164 11854 17220
rect 20300 17164 20860 17220
rect 20916 17164 20926 17220
rect 24994 17164 25004 17220
rect 25060 17164 30940 17220
rect 30996 17164 31500 17220
rect 31556 17164 31566 17220
rect 33170 17164 33180 17220
rect 33236 17164 33740 17220
rect 33796 17164 33806 17220
rect 6738 17052 6748 17108
rect 6804 17052 7420 17108
rect 7476 17052 7486 17108
rect 18834 17052 18844 17108
rect 18900 17052 19404 17108
rect 19460 17052 19852 17108
rect 19908 17052 19918 17108
rect 4050 16940 4060 16996
rect 4116 16940 6860 16996
rect 6916 16940 6926 16996
rect 7074 16940 7084 16996
rect 7140 16940 8988 16996
rect 9044 16940 9054 16996
rect 19852 16884 19908 17052
rect 20300 16996 20356 17164
rect 20066 16940 20076 16996
rect 20132 16940 20356 16996
rect 20524 17052 24668 17108
rect 24724 17052 29148 17108
rect 29204 17052 29214 17108
rect 35410 17052 35420 17108
rect 35476 17052 36428 17108
rect 36484 17052 36494 17108
rect 20524 16884 20580 17052
rect 20738 16940 20748 16996
rect 20804 16940 22540 16996
rect 22596 16940 22606 16996
rect 31714 16940 31724 16996
rect 31780 16940 35532 16996
rect 35588 16940 35598 16996
rect 2482 16828 2492 16884
rect 2548 16828 3388 16884
rect 3444 16828 5740 16884
rect 5796 16828 5806 16884
rect 6066 16828 6076 16884
rect 6132 16828 7868 16884
rect 7924 16828 9772 16884
rect 9828 16828 9838 16884
rect 14018 16828 14028 16884
rect 14084 16828 15036 16884
rect 15092 16828 17500 16884
rect 17556 16828 18508 16884
rect 18564 16828 18574 16884
rect 19852 16828 20580 16884
rect 21858 16828 21868 16884
rect 21924 16828 25452 16884
rect 25508 16828 25518 16884
rect 33394 16828 33404 16884
rect 33460 16828 36428 16884
rect 36484 16828 36494 16884
rect 6178 16716 6188 16772
rect 6244 16716 7420 16772
rect 7476 16716 7756 16772
rect 7812 16716 7822 16772
rect 8194 16716 8204 16772
rect 8260 16716 8764 16772
rect 8820 16716 9324 16772
rect 9380 16716 10668 16772
rect 10724 16716 10734 16772
rect 17042 16716 17052 16772
rect 17108 16716 19068 16772
rect 19124 16716 19134 16772
rect 36306 16716 36316 16772
rect 36372 16716 37772 16772
rect 37828 16716 37838 16772
rect 3500 16604 15148 16660
rect 16146 16604 16156 16660
rect 16212 16604 17388 16660
rect 17444 16604 22204 16660
rect 22260 16604 22270 16660
rect 31602 16604 31612 16660
rect 31668 16604 32732 16660
rect 32788 16604 32798 16660
rect 3500 16548 3556 16604
rect 15092 16548 15148 16604
rect 3490 16492 3500 16548
rect 3556 16492 3566 16548
rect 15092 16492 25228 16548
rect 25284 16492 25294 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 17388 16380 21644 16436
rect 21700 16380 21710 16436
rect 23314 16380 23324 16436
rect 23380 16380 33908 16436
rect 2594 16268 2604 16324
rect 2660 16268 10556 16324
rect 10612 16268 10622 16324
rect 0 16212 800 16240
rect 17388 16212 17444 16380
rect 33852 16324 33908 16380
rect 20178 16268 20188 16324
rect 20244 16268 21308 16324
rect 21364 16268 21374 16324
rect 30146 16268 30156 16324
rect 30212 16268 33628 16324
rect 33684 16268 33694 16324
rect 33852 16268 37100 16324
rect 37156 16268 37166 16324
rect 0 16156 1820 16212
rect 1876 16156 1886 16212
rect 5730 16156 5740 16212
rect 5796 16156 14028 16212
rect 14084 16156 14094 16212
rect 14252 16156 17444 16212
rect 17714 16156 17724 16212
rect 17780 16156 17948 16212
rect 18004 16156 18014 16212
rect 19058 16156 19068 16212
rect 19124 16156 20076 16212
rect 20132 16156 20142 16212
rect 29586 16156 29596 16212
rect 29652 16156 32060 16212
rect 32116 16156 35532 16212
rect 35588 16156 36316 16212
rect 36372 16156 36988 16212
rect 37044 16156 37660 16212
rect 37716 16156 38668 16212
rect 0 16128 800 16156
rect 14252 16100 14308 16156
rect 17724 16100 17780 16156
rect 38612 16100 38668 16156
rect 6962 16044 6972 16100
rect 7028 16044 7868 16100
rect 7924 16044 7934 16100
rect 12898 16044 12908 16100
rect 12964 16044 13244 16100
rect 13300 16044 14308 16100
rect 15092 16044 17780 16100
rect 31154 16044 31164 16100
rect 31220 16044 31500 16100
rect 31556 16044 31566 16100
rect 38612 16044 39900 16100
rect 39956 16044 39966 16100
rect 15092 15988 15148 16044
rect 5954 15932 5964 15988
rect 6020 15932 7084 15988
rect 7140 15932 7150 15988
rect 8082 15932 8092 15988
rect 8148 15932 8652 15988
rect 8708 15932 15148 15988
rect 15362 15932 15372 15988
rect 15428 15932 16940 15988
rect 16996 15932 17006 15988
rect 18946 15932 18956 15988
rect 19012 15932 19740 15988
rect 19796 15932 21420 15988
rect 21476 15932 21980 15988
rect 22036 15932 22046 15988
rect 30930 15932 30940 15988
rect 30996 15932 31388 15988
rect 31444 15932 33068 15988
rect 33124 15932 33134 15988
rect 7186 15820 7196 15876
rect 7252 15820 7644 15876
rect 7700 15820 7710 15876
rect 13122 15820 13132 15876
rect 13188 15820 13468 15876
rect 13524 15820 14252 15876
rect 14308 15820 14700 15876
rect 14756 15820 14766 15876
rect 30706 15820 30716 15876
rect 30772 15820 31164 15876
rect 31220 15820 31230 15876
rect 31378 15820 31388 15876
rect 31444 15820 34860 15876
rect 34916 15820 34926 15876
rect 35970 15820 35980 15876
rect 36036 15820 37212 15876
rect 37268 15820 38668 15876
rect 38724 15820 39228 15876
rect 39284 15820 39294 15876
rect 28812 15708 29932 15764
rect 29988 15708 29998 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 12450 15596 12460 15652
rect 12516 15596 15260 15652
rect 15316 15596 15326 15652
rect 25218 15596 25228 15652
rect 25284 15596 26012 15652
rect 26068 15596 26796 15652
rect 26852 15596 27804 15652
rect 27860 15596 27870 15652
rect 28812 15540 28868 15708
rect 6178 15484 6188 15540
rect 6244 15484 6860 15540
rect 6916 15484 6926 15540
rect 7746 15484 7756 15540
rect 7812 15484 9548 15540
rect 9604 15484 9614 15540
rect 9986 15484 9996 15540
rect 10052 15484 12796 15540
rect 12852 15484 14924 15540
rect 14980 15484 14990 15540
rect 15820 15484 28868 15540
rect 28924 15596 32396 15652
rect 32452 15596 32462 15652
rect 3154 15372 3164 15428
rect 3220 15372 6748 15428
rect 6804 15372 6814 15428
rect 14578 15372 14588 15428
rect 14644 15372 15596 15428
rect 15652 15372 15662 15428
rect 15820 15316 15876 15484
rect 28924 15428 28980 15596
rect 30258 15484 30268 15540
rect 30324 15484 31724 15540
rect 31780 15484 33180 15540
rect 33236 15484 33246 15540
rect 21606 15372 21644 15428
rect 21700 15372 21710 15428
rect 22082 15372 22092 15428
rect 22148 15372 22708 15428
rect 22652 15316 22708 15372
rect 26852 15372 28980 15428
rect 35746 15372 35756 15428
rect 35812 15372 37100 15428
rect 37156 15372 37166 15428
rect 26852 15316 26908 15372
rect 11778 15260 11788 15316
rect 11844 15260 15876 15316
rect 19954 15260 19964 15316
rect 20020 15260 20972 15316
rect 21028 15260 21038 15316
rect 21410 15260 21420 15316
rect 21476 15260 22316 15316
rect 22372 15260 22382 15316
rect 22642 15260 22652 15316
rect 22708 15260 26908 15316
rect 28018 15260 28028 15316
rect 28084 15260 28588 15316
rect 28644 15260 35868 15316
rect 35924 15260 35934 15316
rect 5282 15148 5292 15204
rect 5348 15148 6300 15204
rect 6356 15148 6366 15204
rect 10322 15148 10332 15204
rect 10388 15148 10892 15204
rect 10948 15148 19404 15204
rect 19460 15148 20076 15204
rect 20132 15148 26460 15204
rect 26516 15148 26526 15204
rect 27906 15148 27916 15204
rect 27972 15148 29260 15204
rect 29316 15148 30156 15204
rect 30212 15148 30222 15204
rect 14466 14924 14476 14980
rect 14532 14924 22092 14980
rect 22148 14924 22158 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 21186 14812 21196 14868
rect 21252 14812 24220 14868
rect 24276 14812 24286 14868
rect 19842 14700 19852 14756
rect 19908 14700 21644 14756
rect 21700 14700 21710 14756
rect 0 14644 800 14672
rect 0 14588 1708 14644
rect 1764 14588 1774 14644
rect 12002 14588 12012 14644
rect 12068 14588 12460 14644
rect 12516 14588 27132 14644
rect 27188 14588 27198 14644
rect 0 14560 800 14588
rect 5506 14476 5516 14532
rect 5572 14476 16156 14532
rect 16212 14476 16222 14532
rect 16370 14476 16380 14532
rect 16436 14476 19068 14532
rect 19124 14476 21644 14532
rect 21700 14476 21868 14532
rect 21924 14476 21934 14532
rect 28914 14476 28924 14532
rect 28980 14476 30156 14532
rect 30212 14476 33292 14532
rect 33348 14476 33358 14532
rect 16380 14420 16436 14476
rect 15250 14364 15260 14420
rect 15316 14364 16436 14420
rect 20066 14364 20076 14420
rect 20132 14364 20412 14420
rect 20468 14364 20478 14420
rect 13906 14252 13916 14308
rect 13972 14252 14252 14308
rect 14308 14252 14318 14308
rect 19954 14252 19964 14308
rect 20020 14252 20972 14308
rect 21028 14252 21252 14308
rect 21410 14252 21420 14308
rect 21476 14252 22540 14308
rect 22596 14252 22606 14308
rect 25666 14252 25676 14308
rect 25732 14252 26684 14308
rect 26740 14252 28588 14308
rect 28644 14252 30716 14308
rect 30772 14252 30782 14308
rect 35858 14252 35868 14308
rect 35924 14252 47852 14308
rect 47908 14252 47918 14308
rect 21196 14196 21252 14252
rect 49200 14196 50000 14224
rect 2258 14140 2268 14196
rect 2324 14140 8428 14196
rect 8484 14140 8494 14196
rect 9874 14140 9884 14196
rect 9940 14140 10780 14196
rect 10836 14140 11228 14196
rect 11284 14140 15932 14196
rect 15988 14140 16492 14196
rect 16548 14140 16558 14196
rect 21196 14140 26460 14196
rect 26516 14140 27244 14196
rect 27300 14140 27580 14196
rect 27636 14140 27646 14196
rect 47618 14140 47628 14196
rect 47684 14140 48188 14196
rect 48244 14140 50000 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 49200 14112 50000 14140
rect 21522 13916 21532 13972
rect 21588 13916 28924 13972
rect 28980 13916 28990 13972
rect 27906 13804 27916 13860
rect 27972 13804 28476 13860
rect 28532 13804 28542 13860
rect 30818 13804 30828 13860
rect 30884 13804 31612 13860
rect 31668 13804 31678 13860
rect 2258 13692 2268 13748
rect 2324 13692 3500 13748
rect 3556 13692 3566 13748
rect 20514 13692 20524 13748
rect 20580 13692 20860 13748
rect 20916 13692 23604 13748
rect 23548 13636 23604 13692
rect 8194 13580 8204 13636
rect 8260 13580 9660 13636
rect 9716 13580 9726 13636
rect 20290 13580 20300 13636
rect 20356 13580 21532 13636
rect 21588 13580 21756 13636
rect 21812 13580 21822 13636
rect 23538 13580 23548 13636
rect 23604 13580 24668 13636
rect 24724 13580 24734 13636
rect 26338 13468 26348 13524
rect 26404 13468 29708 13524
rect 29764 13468 29774 13524
rect 31350 13468 31388 13524
rect 31444 13468 31454 13524
rect 27804 13412 27860 13468
rect 21718 13356 21756 13412
rect 21812 13356 21822 13412
rect 27794 13356 27804 13412
rect 27860 13356 27870 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 30594 13244 30604 13300
rect 30660 13244 31052 13300
rect 31108 13244 31118 13300
rect 0 13076 800 13104
rect 0 13020 1820 13076
rect 1876 13020 1886 13076
rect 17378 13020 17388 13076
rect 17444 13020 20300 13076
rect 20356 13020 20366 13076
rect 28578 13020 28588 13076
rect 28644 13020 29372 13076
rect 29428 13020 29438 13076
rect 31266 13020 31276 13076
rect 31332 13020 32732 13076
rect 32788 13020 32798 13076
rect 34178 13020 34188 13076
rect 34244 13020 34860 13076
rect 34916 13020 34926 13076
rect 0 12992 800 13020
rect 10434 12908 10444 12964
rect 10500 12908 11452 12964
rect 11508 12908 11518 12964
rect 12674 12908 12684 12964
rect 12740 12908 14588 12964
rect 14644 12908 14654 12964
rect 16706 12908 16716 12964
rect 16772 12908 21532 12964
rect 21588 12908 21598 12964
rect 30034 12908 30044 12964
rect 30100 12908 30268 12964
rect 30324 12908 30334 12964
rect 27234 12796 27244 12852
rect 27300 12796 27692 12852
rect 27748 12796 27758 12852
rect 34188 12740 34244 13020
rect 23650 12684 23660 12740
rect 23716 12684 30492 12740
rect 30548 12684 31500 12740
rect 31556 12684 34244 12740
rect 30034 12572 30044 12628
rect 30100 12572 31052 12628
rect 31108 12572 31118 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 11666 12348 11676 12404
rect 11732 12348 12124 12404
rect 12180 12348 14140 12404
rect 14196 12348 14206 12404
rect 11442 12236 11452 12292
rect 11508 12236 13356 12292
rect 13412 12236 13916 12292
rect 13972 12236 13982 12292
rect 20514 12236 20524 12292
rect 20580 12236 21420 12292
rect 21476 12236 21486 12292
rect 27346 12124 27356 12180
rect 27412 12124 27916 12180
rect 27972 12124 28588 12180
rect 28644 12124 29260 12180
rect 29316 12124 30380 12180
rect 30436 12124 30446 12180
rect 2258 12012 2268 12068
rect 2324 12012 8428 12068
rect 18050 12012 18060 12068
rect 18116 12012 19180 12068
rect 19236 12012 19246 12068
rect 20962 12012 20972 12068
rect 21028 12012 23772 12068
rect 23828 12012 23838 12068
rect 8372 11956 8428 12012
rect 20972 11956 21028 12012
rect 8372 11900 21028 11956
rect 30146 11900 30156 11956
rect 30212 11900 32228 11956
rect 23538 11788 23548 11844
rect 23604 11788 25452 11844
rect 25508 11788 26348 11844
rect 26404 11788 26796 11844
rect 26852 11788 29204 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 29148 11732 29204 11788
rect 31892 11732 31948 11844
rect 32004 11788 32014 11844
rect 6066 11676 6076 11732
rect 6132 11676 9772 11732
rect 9828 11676 15148 11732
rect 15204 11676 15484 11732
rect 15540 11676 15550 11732
rect 29138 11676 29148 11732
rect 29204 11676 30940 11732
rect 30996 11676 31948 11732
rect 32172 11732 32228 11900
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 32172 11676 33964 11732
rect 34020 11676 34030 11732
rect 11554 11564 11564 11620
rect 11620 11564 12796 11620
rect 12852 11564 14812 11620
rect 14868 11564 15820 11620
rect 15876 11564 15886 11620
rect 0 11508 800 11536
rect 0 11452 1820 11508
rect 1876 11452 1886 11508
rect 2370 11452 2380 11508
rect 2436 11452 15148 11508
rect 15586 11452 15596 11508
rect 15652 11452 16492 11508
rect 16548 11452 23660 11508
rect 23716 11452 23726 11508
rect 30594 11452 30604 11508
rect 30660 11452 31612 11508
rect 31668 11452 31678 11508
rect 0 11424 800 11452
rect 15092 11396 15148 11452
rect 15092 11340 20748 11396
rect 20804 11340 21868 11396
rect 21924 11340 25676 11396
rect 25732 11340 25742 11396
rect 32172 11172 32228 11676
rect 9426 11116 9436 11172
rect 9492 11116 11788 11172
rect 11844 11116 11854 11172
rect 26898 11116 26908 11172
rect 26964 11116 32228 11172
rect 32722 11116 32732 11172
rect 32788 11116 34524 11172
rect 34580 11116 34590 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 15810 10780 15820 10836
rect 15876 10780 16492 10836
rect 16548 10780 26236 10836
rect 26292 10780 27244 10836
rect 27300 10780 27310 10836
rect 2258 10668 2268 10724
rect 2324 10668 3052 10724
rect 3108 10668 15148 10724
rect 19394 10668 19404 10724
rect 19460 10668 20076 10724
rect 20132 10668 20142 10724
rect 15092 10612 15148 10668
rect 15092 10556 20244 10612
rect 12002 10332 12012 10388
rect 12068 10332 15372 10388
rect 15428 10332 15438 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 20188 10164 20244 10556
rect 29138 10444 29148 10500
rect 29204 10444 29708 10500
rect 29764 10444 32732 10500
rect 32788 10444 32798 10500
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 20178 10108 20188 10164
rect 20244 10108 25004 10164
rect 25060 10108 25070 10164
rect 12450 9996 12460 10052
rect 12516 9996 20972 10052
rect 21028 9996 21038 10052
rect 22418 9996 22428 10052
rect 22484 9996 23100 10052
rect 23156 9996 23166 10052
rect 26898 9996 26908 10052
rect 26964 9996 26974 10052
rect 0 9940 800 9968
rect 26908 9940 26964 9996
rect 0 9884 1820 9940
rect 1876 9884 1886 9940
rect 11666 9884 11676 9940
rect 11732 9884 12124 9940
rect 12180 9884 12190 9940
rect 14130 9884 14140 9940
rect 14196 9884 15372 9940
rect 15428 9884 26964 9940
rect 0 9856 800 9884
rect 8754 9772 8764 9828
rect 8820 9772 9660 9828
rect 9716 9772 9726 9828
rect 14354 9772 14364 9828
rect 14420 9772 15708 9828
rect 15764 9772 15774 9828
rect 20066 9772 20076 9828
rect 20132 9772 20524 9828
rect 20580 9772 21868 9828
rect 21924 9772 21934 9828
rect 22194 9772 22204 9828
rect 22260 9772 22764 9828
rect 22820 9772 23548 9828
rect 23604 9772 24332 9828
rect 24388 9772 24398 9828
rect 9874 9660 9884 9716
rect 9940 9660 17388 9716
rect 17444 9660 18620 9716
rect 18676 9660 20188 9716
rect 20244 9660 20254 9716
rect 24434 9660 24444 9716
rect 24500 9660 25900 9716
rect 25956 9660 25966 9716
rect 20066 9548 20076 9604
rect 20132 9548 20188 9604
rect 20244 9548 20254 9604
rect 20962 9548 20972 9604
rect 21028 9548 30268 9604
rect 30324 9548 32172 9604
rect 32228 9548 32238 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 2034 9212 2044 9268
rect 2100 9212 5516 9268
rect 5572 9212 5582 9268
rect 9650 9212 9660 9268
rect 9716 9212 11788 9268
rect 11844 9212 12684 9268
rect 12740 9212 14812 9268
rect 14868 9212 15932 9268
rect 15988 9212 16940 9268
rect 16996 9212 17006 9268
rect 20738 9100 20748 9156
rect 20804 9100 22204 9156
rect 22260 9100 22270 9156
rect 32274 9100 32284 9156
rect 32340 9100 47852 9156
rect 47908 9100 47918 9156
rect 19730 8988 19740 9044
rect 19796 8988 20524 9044
rect 20580 8988 20590 9044
rect 21298 8988 21308 9044
rect 21364 8988 21868 9044
rect 21924 8988 21934 9044
rect 21308 8932 21364 8988
rect 19170 8876 19180 8932
rect 19236 8876 20076 8932
rect 20132 8876 21364 8932
rect 26226 8876 26236 8932
rect 26292 8876 27132 8932
rect 27188 8876 35980 8932
rect 36036 8876 36046 8932
rect 49200 8820 50000 8848
rect 47618 8764 47628 8820
rect 47684 8764 48188 8820
rect 48244 8764 50000 8820
rect 49200 8736 50000 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 0 8372 800 8400
rect 0 8316 1708 8372
rect 1764 8316 2492 8372
rect 2548 8316 2558 8372
rect 22642 8316 22652 8372
rect 22708 8316 23660 8372
rect 23716 8316 23726 8372
rect 0 8288 800 8316
rect 22978 8204 22988 8260
rect 23044 8204 26348 8260
rect 26404 8204 26414 8260
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 21074 7644 21084 7700
rect 21140 7644 21868 7700
rect 21924 7644 31164 7700
rect 31220 7644 31230 7700
rect 1698 7308 1708 7364
rect 1764 7308 2492 7364
rect 2548 7308 2558 7364
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 0 6804 800 6832
rect 0 6748 1708 6804
rect 1764 6748 1774 6804
rect 0 6720 800 6748
rect 16818 6636 16828 6692
rect 16884 6636 20188 6692
rect 20244 6636 20254 6692
rect 23650 6636 23660 6692
rect 23716 6636 24220 6692
rect 24276 6636 28700 6692
rect 28756 6636 28766 6692
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 28242 5964 28252 6020
rect 28308 5964 29036 6020
rect 29092 5964 29102 6020
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 0 5236 800 5264
rect 0 5180 1820 5236
rect 1876 5180 1886 5236
rect 22642 5180 22652 5236
rect 22708 5180 24108 5236
rect 24164 5180 24174 5236
rect 0 5152 800 5180
rect 35970 4956 35980 5012
rect 36036 4956 37436 5012
rect 37492 4956 37502 5012
rect 39778 4956 39788 5012
rect 39844 4956 42028 5012
rect 42084 4956 42094 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 40338 4508 40348 4564
rect 40404 4508 41244 4564
rect 41300 4508 41310 4564
rect 44482 4508 44492 4564
rect 44548 4508 47852 4564
rect 47908 4508 47918 4564
rect 1698 4172 1708 4228
rect 1764 4172 2492 4228
rect 2548 4172 2558 4228
rect 8754 4060 8764 4116
rect 8820 4060 9772 4116
rect 9828 4060 9838 4116
rect 12786 4060 12796 4116
rect 12852 4060 14028 4116
rect 14084 4060 14094 4116
rect 26898 4060 26908 4116
rect 26964 4060 28140 4116
rect 28196 4060 28206 4116
rect 32946 4060 32956 4116
rect 33012 4060 34188 4116
rect 34244 4060 34254 4116
rect 41010 4060 41020 4116
rect 41076 4060 42252 4116
rect 42308 4060 42318 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 0 3668 800 3696
rect 0 3612 1708 3668
rect 1764 3612 1774 3668
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 38994 3612 39004 3668
rect 39060 3612 40012 3668
rect 40068 3612 40078 3668
rect 42018 3612 42028 3668
rect 42084 3612 42812 3668
rect 42868 3612 42878 3668
rect 46274 3612 46284 3668
rect 46340 3612 47852 3668
rect 47908 3612 47918 3668
rect 0 3584 800 3612
rect 17826 3500 17836 3556
rect 17892 3500 19180 3556
rect 19236 3500 20076 3556
rect 20132 3500 20142 3556
rect 26114 3500 26124 3556
rect 26180 3500 27244 3556
rect 27300 3500 28476 3556
rect 28532 3500 28542 3556
rect 32610 3500 32620 3556
rect 32676 3500 33628 3556
rect 33684 3500 33694 3556
rect 43474 3500 43484 3556
rect 43540 3500 45724 3556
rect 45780 3500 46620 3556
rect 46676 3500 46686 3556
rect 49200 3444 50000 3472
rect 28914 3388 28924 3444
rect 28980 3388 30044 3444
rect 30100 3388 30110 3444
rect 30930 3388 30940 3444
rect 30996 3388 33740 3444
rect 33796 3388 33806 3444
rect 35522 3388 35532 3444
rect 35588 3388 36204 3444
rect 36260 3388 36270 3444
rect 48178 3388 48188 3444
rect 48244 3388 50000 3444
rect 49200 3360 50000 3388
rect 1698 3276 1708 3332
rect 1764 3276 2940 3332
rect 2996 3276 3006 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 0 2100 800 2128
rect 0 2044 1708 2100
rect 1764 2044 1774 2100
rect 0 2016 800 2044
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 12236 45052 12292 45108
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 27468 44380 27524 44436
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 18060 42924 18116 42980
rect 18060 42476 18116 42532
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 27692 42028 27748 42084
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 27468 38556 27524 38612
rect 27692 38556 27748 38612
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 4956 38108 5012 38164
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 13916 37324 13972 37380
rect 9772 37100 9828 37156
rect 4956 36876 5012 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 14028 36540 14084 36596
rect 13916 36204 13972 36260
rect 12236 36092 12292 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 19628 35868 19684 35924
rect 14028 35644 14084 35700
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 10780 35084 10836 35140
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 22876 33404 22932 33460
rect 9996 33292 10052 33348
rect 9772 33180 9828 33236
rect 19404 32956 19460 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 26908 32844 26964 32900
rect 10780 32620 10836 32676
rect 34412 32732 34468 32788
rect 9212 32284 9268 32340
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 34188 32060 34244 32116
rect 8316 31500 8372 31556
rect 8540 31500 8596 31556
rect 26908 31388 26964 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 8764 31276 8820 31332
rect 14252 30828 14308 30884
rect 8204 30716 8260 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 34188 30492 34244 30548
rect 14252 30380 14308 30436
rect 33628 30380 33684 30436
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 19404 29148 19460 29204
rect 19628 29148 19684 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 8764 28476 8820 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 8540 27804 8596 27860
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19292 26908 19348 26964
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 9212 26012 9268 26068
rect 9996 26012 10052 26068
rect 22876 26012 22932 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 8316 25116 8372 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 14252 25004 14308 25060
rect 19292 25004 19348 25060
rect 34300 25004 34356 25060
rect 8204 24780 8260 24836
rect 33628 24444 33684 24500
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 34412 24220 34468 24276
rect 34300 24108 34356 24164
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 15596 22428 15652 22484
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 21756 21868 21812 21924
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 14140 21084 14196 21140
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 15596 20076 15652 20132
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 31388 18956 31444 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 15596 18620 15652 18676
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 31388 15820 31444 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 21644 15372 21700 15428
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 21644 14476 21700 14532
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 31388 13468 31444 13524
rect 21756 13356 21812 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 14140 12348 14196 12404
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 20188 10108 20244 10164
rect 20972 9996 21028 10052
rect 20188 9548 20244 9604
rect 20972 9548 21028 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 12236 45108 12292 45118
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4956 38164 5012 38174
rect 4956 36932 5012 38108
rect 4956 36866 5012 36876
rect 9772 37156 9828 37166
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 9772 33236 9828 37100
rect 12236 36148 12292 45052
rect 19808 43932 20128 45444
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 18060 42980 18116 42990
rect 18060 42532 18116 42924
rect 18060 42466 18116 42476
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 27468 44436 27524 44446
rect 27468 38612 27524 44380
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 27468 38546 27524 38556
rect 27692 42084 27748 42094
rect 27692 38612 27748 42028
rect 27692 38546 27748 38556
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 13916 37380 13972 37390
rect 13916 36260 13972 37324
rect 13916 36194 13972 36204
rect 14028 36596 14084 36606
rect 12236 36082 12292 36092
rect 14028 35700 14084 36540
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 14028 35634 14084 35644
rect 19628 35924 19684 35934
rect 10780 35140 10836 35150
rect 9772 33170 9828 33180
rect 9996 33348 10052 33358
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 9212 32340 9268 32350
rect 8316 31556 8372 31566
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 8204 30772 8260 30782
rect 8204 24836 8260 30716
rect 8316 25172 8372 31500
rect 8540 31556 8596 31566
rect 8540 27860 8596 31500
rect 8764 31332 8820 31342
rect 8764 28532 8820 31276
rect 8764 28466 8820 28476
rect 8540 27794 8596 27804
rect 9212 26068 9268 32284
rect 9212 26002 9268 26012
rect 9996 26068 10052 33292
rect 10780 32676 10836 35084
rect 10780 32610 10836 32620
rect 19404 33012 19460 33022
rect 9996 26002 10052 26012
rect 14252 30884 14308 30894
rect 14252 30436 14308 30828
rect 8316 25106 8372 25116
rect 14252 25060 14308 30380
rect 19404 29204 19460 32956
rect 19404 29138 19460 29148
rect 19628 29204 19684 35868
rect 19628 29138 19684 29148
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 14252 24994 14308 25004
rect 19292 26964 19348 26974
rect 19292 25060 19348 26908
rect 19292 24994 19348 25004
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 22876 33460 22932 33470
rect 22876 26068 22932 33404
rect 26908 32900 26964 32910
rect 26908 31444 26964 32844
rect 34412 32788 34468 32798
rect 26908 31378 26964 31388
rect 34188 32116 34244 32126
rect 34188 30548 34244 32060
rect 34188 30482 34244 30492
rect 22876 26002 22932 26012
rect 33628 30436 33684 30446
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 8204 24770 8260 24780
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 23548 20128 25060
rect 33628 24500 33684 30380
rect 33628 24434 33684 24444
rect 34300 25060 34356 25070
rect 34300 24164 34356 25004
rect 34412 24276 34468 32732
rect 34412 24210 34468 24220
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 34300 24098 34356 24108
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 15596 22484 15652 22494
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 14140 21140 14196 21150
rect 14140 12404 14196 21084
rect 15596 20132 15652 22428
rect 15596 18676 15652 20076
rect 15596 18610 15652 18620
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 14140 12338 14196 12348
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 21756 21924 21812 21934
rect 21644 15428 21700 15438
rect 21644 14532 21700 15372
rect 21644 14466 21700 14476
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 21756 13412 21812 21868
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 31388 19012 31444 19022
rect 31388 15876 31444 18956
rect 31388 13524 31444 15820
rect 31388 13458 31444 13468
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 21756 13346 21812 13356
rect 35168 13356 35488 14868
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 20188 10164 20244 10174
rect 20188 9604 20244 10108
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 20188 9538 20244 9548
rect 20972 10052 21028 10062
rect 20972 9604 21028 9996
rect 20972 9538 21028 9548
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _400_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _401_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20272 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _402_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _403_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18928 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1698431365
transform 1 0 23632 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _405_
timestamp 1698431365
transform 1 0 22624 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _406_
timestamp 1698431365
transform 1 0 23632 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _407_
timestamp 1698431365
transform 1 0 25424 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _408_
timestamp 1698431365
transform -1 0 29120 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_
timestamp 1698431365
transform -1 0 29680 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _410_
timestamp 1698431365
transform 1 0 30128 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _411_
timestamp 1698431365
transform -1 0 30464 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _412_
timestamp 1698431365
transform -1 0 34608 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _413_
timestamp 1698431365
transform 1 0 31360 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _414_
timestamp 1698431365
transform 1 0 33712 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _415_
timestamp 1698431365
transform 1 0 33936 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _416_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _417_
timestamp 1698431365
transform 1 0 24192 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _418_
timestamp 1698431365
transform 1 0 32592 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _419_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6944 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _420_
timestamp 1698431365
transform -1 0 16240 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _421_
timestamp 1698431365
transform -1 0 12880 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _422_
timestamp 1698431365
transform -1 0 14560 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _423_
timestamp 1698431365
transform 1 0 15008 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _424_
timestamp 1698431365
transform 1 0 7280 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _425_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7616 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _426_
timestamp 1698431365
transform -1 0 21616 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _427_
timestamp 1698431365
transform 1 0 30016 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _428_
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _429_
timestamp 1698431365
transform -1 0 36176 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _430_
timestamp 1698431365
transform 1 0 35168 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _431_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28000 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _432_
timestamp 1698431365
transform 1 0 26656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _433_
timestamp 1698431365
transform 1 0 27664 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _434_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _435_
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _436_
timestamp 1698431365
transform 1 0 33264 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _437_
timestamp 1698431365
transform -1 0 40432 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _438_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39312 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _439_
timestamp 1698431365
transform -1 0 41888 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _440_
timestamp 1698431365
transform 1 0 40768 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _441_
timestamp 1698431365
transform -1 0 42224 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _442_
timestamp 1698431365
transform 1 0 42672 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _443_
timestamp 1698431365
transform -1 0 43792 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _444_
timestamp 1698431365
transform 1 0 43344 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _445_
timestamp 1698431365
transform 1 0 20496 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _446_
timestamp 1698431365
transform 1 0 25760 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _447_
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _448_
timestamp 1698431365
transform 1 0 29344 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _449_
timestamp 1698431365
transform 1 0 31584 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _450_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6496 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _451_
timestamp 1698431365
transform -1 0 8400 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _452_
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _453_
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _454_
timestamp 1698431365
transform -1 0 22960 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _455_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23856 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _456_
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _457_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _458_
timestamp 1698431365
transform 1 0 28896 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _459_
timestamp 1698431365
transform 1 0 31136 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _460_
timestamp 1698431365
transform 1 0 19040 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _461_
timestamp 1698431365
transform 1 0 44800 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _462_
timestamp 1698431365
transform -1 0 11312 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _463_
timestamp 1698431365
transform -1 0 10640 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _464_
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _465_
timestamp 1698431365
transform 1 0 15792 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _466_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38976 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _467_
timestamp 1698431365
transform -1 0 21280 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _468_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12880 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _469_
timestamp 1698431365
transform -1 0 11200 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _470_
timestamp 1698431365
transform -1 0 9296 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _471_
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _472_
timestamp 1698431365
transform 1 0 9968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _473_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _474_
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _475_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11760 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _476_
timestamp 1698431365
transform 1 0 13664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _477_
timestamp 1698431365
transform 1 0 19040 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _478_
timestamp 1698431365
transform 1 0 8512 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12880 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _480_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _481_
timestamp 1698431365
transform 1 0 11536 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _482_
timestamp 1698431365
transform 1 0 10864 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _483_
timestamp 1698431365
transform 1 0 11312 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _484_
timestamp 1698431365
transform 1 0 9296 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _485_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13776 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _486_
timestamp 1698431365
transform 1 0 19712 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _487_
timestamp 1698431365
transform 1 0 10416 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _488_
timestamp 1698431365
transform -1 0 16576 0 -1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _489_
timestamp 1698431365
transform 1 0 13664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _490_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _491_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11536 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _492_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12656 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _493_
timestamp 1698431365
transform -1 0 16912 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _494_
timestamp 1698431365
transform 1 0 19936 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _495_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20160 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _496_
timestamp 1698431365
transform 1 0 8288 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _497_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _498_
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _499_
timestamp 1698431365
transform 1 0 10528 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _500_
timestamp 1698431365
transform 1 0 13664 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _501_
timestamp 1698431365
transform 1 0 14448 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _502_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _503_
timestamp 1698431365
transform 1 0 11760 0 -1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _504_
timestamp 1698431365
transform 1 0 14896 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _505_
timestamp 1698431365
transform -1 0 16352 0 -1 37632
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _506_
timestamp 1698431365
transform 1 0 12656 0 -1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _507_
timestamp 1698431365
transform 1 0 10192 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _508_
timestamp 1698431365
transform 1 0 12208 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _509_
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _510_
timestamp 1698431365
transform 1 0 12768 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _511_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _512_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15792 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _513_
timestamp 1698431365
transform -1 0 10304 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _514_
timestamp 1698431365
transform -1 0 8288 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _515_
timestamp 1698431365
transform 1 0 5600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _516_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12656 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _517_
timestamp 1698431365
transform 1 0 8624 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _518_
timestamp 1698431365
transform -1 0 9072 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _519_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _520_
timestamp 1698431365
transform 1 0 11424 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _521_
timestamp 1698431365
transform -1 0 18704 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _522_
timestamp 1698431365
transform 1 0 17808 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _523_
timestamp 1698431365
transform -1 0 20160 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _524_
timestamp 1698431365
transform -1 0 14448 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _525_
timestamp 1698431365
transform -1 0 8176 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _526_
timestamp 1698431365
transform 1 0 6608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _527_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14560 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _528_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _529_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17808 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _530_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18368 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _531_
timestamp 1698431365
transform 1 0 15904 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _532_
timestamp 1698431365
transform -1 0 10080 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _533_
timestamp 1698431365
transform -1 0 12992 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _534_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _535_
timestamp 1698431365
transform 1 0 18704 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _536_
timestamp 1698431365
transform 1 0 9296 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _537_
timestamp 1698431365
transform -1 0 9296 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _538_
timestamp 1698431365
transform -1 0 10640 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _539_
timestamp 1698431365
transform -1 0 9072 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _540_
timestamp 1698431365
transform -1 0 9968 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _541_
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _542_
timestamp 1698431365
transform 1 0 16128 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _543_
timestamp 1698431365
transform 1 0 15120 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _544_
timestamp 1698431365
transform 1 0 16912 0 1 26656
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _545_
timestamp 1698431365
transform 1 0 15904 0 1 36064
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _546_
timestamp 1698431365
transform 1 0 12096 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _547_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8960 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _548_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9968 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _549_
timestamp 1698431365
transform -1 0 9184 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _550_
timestamp 1698431365
transform 1 0 7504 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _551_
timestamp 1698431365
transform -1 0 24640 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _552_
timestamp 1698431365
transform 1 0 14560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _553_
timestamp 1698431365
transform 1 0 15904 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _554_
timestamp 1698431365
transform 1 0 14336 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _555_
timestamp 1698431365
transform -1 0 12992 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _556_
timestamp 1698431365
transform 1 0 18256 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _557_
timestamp 1698431365
transform -1 0 12768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _558_
timestamp 1698431365
transform -1 0 10640 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _559_
timestamp 1698431365
transform 1 0 7392 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _560_
timestamp 1698431365
transform -1 0 20048 0 -1 28224
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _561_
timestamp 1698431365
transform -1 0 12768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _562_
timestamp 1698431365
transform -1 0 14336 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _563_
timestamp 1698431365
transform 1 0 9856 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _564_
timestamp 1698431365
transform 1 0 17248 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _565_
timestamp 1698431365
transform -1 0 12768 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _566_
timestamp 1698431365
transform -1 0 9968 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _567_
timestamp 1698431365
transform 1 0 7504 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _568_
timestamp 1698431365
transform 1 0 14112 0 -1 28224
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _569_
timestamp 1698431365
transform -1 0 17024 0 -1 39200
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _570_
timestamp 1698431365
transform -1 0 19712 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _571_
timestamp 1698431365
transform -1 0 19712 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _572_
timestamp 1698431365
transform -1 0 18592 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _573_
timestamp 1698431365
transform -1 0 10640 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _574_
timestamp 1698431365
transform 1 0 5600 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _575_
timestamp 1698431365
transform -1 0 15456 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _576_
timestamp 1698431365
transform 1 0 11312 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _577_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15568 0 -1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _578_
timestamp 1698431365
transform 1 0 14448 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _579_
timestamp 1698431365
transform -1 0 10416 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _580_
timestamp 1698431365
transform 1 0 14448 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _581_
timestamp 1698431365
transform -1 0 22512 0 -1 31360
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _582_
timestamp 1698431365
transform -1 0 12432 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _583_
timestamp 1698431365
transform -1 0 9184 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _584_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _585_
timestamp 1698431365
transform 1 0 22176 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _586_
timestamp 1698431365
transform -1 0 23408 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _587_
timestamp 1698431365
transform 1 0 22960 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _588_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33824 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _589_
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _590_
timestamp 1698431365
transform 1 0 34608 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _591_
timestamp 1698431365
transform 1 0 34608 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _592_
timestamp 1698431365
transform 1 0 36176 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _593_
timestamp 1698431365
transform 1 0 28896 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _594_
timestamp 1698431365
transform 1 0 33824 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _595_
timestamp 1698431365
transform 1 0 31360 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _596_
timestamp 1698431365
transform 1 0 34608 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _597_
timestamp 1698431365
transform -1 0 36064 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _598_
timestamp 1698431365
transform 1 0 36400 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _599_
timestamp 1698431365
transform 1 0 23072 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _600_
timestamp 1698431365
transform 1 0 34272 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _601_
timestamp 1698431365
transform 1 0 39760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _602_
timestamp 1698431365
transform 1 0 38864 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _603_
timestamp 1698431365
transform 1 0 39312 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _604_
timestamp 1698431365
transform 1 0 17248 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _605_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _606_
timestamp 1698431365
transform -1 0 20160 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _607_
timestamp 1698431365
transform -1 0 16128 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _608_
timestamp 1698431365
transform -1 0 13552 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _609_
timestamp 1698431365
transform -1 0 8736 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _610_
timestamp 1698431365
transform 1 0 23408 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _611_
timestamp 1698431365
transform -1 0 10080 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _612_
timestamp 1698431365
transform -1 0 6160 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _613_
timestamp 1698431365
transform -1 0 5152 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _614_
timestamp 1698431365
transform 1 0 4704 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _615_
timestamp 1698431365
transform -1 0 10752 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _616_
timestamp 1698431365
transform 1 0 6608 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _617_
timestamp 1698431365
transform -1 0 4704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _618_
timestamp 1698431365
transform -1 0 3136 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _619_
timestamp 1698431365
transform 1 0 10640 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _620_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4256 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _621_
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _622_
timestamp 1698431365
transform -1 0 9184 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _623_
timestamp 1698431365
transform -1 0 8624 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _624_
timestamp 1698431365
transform -1 0 8960 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _625_
timestamp 1698431365
transform -1 0 7728 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _626_
timestamp 1698431365
transform -1 0 5264 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _627_
timestamp 1698431365
transform -1 0 4256 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _628_
timestamp 1698431365
transform 1 0 3136 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _629_
timestamp 1698431365
transform 1 0 26544 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _630_
timestamp 1698431365
transform -1 0 12208 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _631_
timestamp 1698431365
transform 1 0 9744 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _632_
timestamp 1698431365
transform 1 0 10304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _633_
timestamp 1698431365
transform 1 0 2688 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _634_
timestamp 1698431365
transform 1 0 4256 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _635_
timestamp 1698431365
transform 1 0 34272 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _636_
timestamp 1698431365
transform -1 0 24528 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _637_
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _638_
timestamp 1698431365
transform -1 0 26432 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _639_
timestamp 1698431365
transform -1 0 12768 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _640_
timestamp 1698431365
transform 1 0 10304 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _641_
timestamp 1698431365
transform -1 0 12096 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _642_
timestamp 1698431365
transform 1 0 20608 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _643_
timestamp 1698431365
transform -1 0 14112 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _644_
timestamp 1698431365
transform -1 0 8400 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _645_
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _646_
timestamp 1698431365
transform -1 0 10080 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _647_
timestamp 1698431365
transform 1 0 7728 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _648_
timestamp 1698431365
transform -1 0 22736 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _649_
timestamp 1698431365
transform -1 0 16352 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _650_
timestamp 1698431365
transform -1 0 11200 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _651_
timestamp 1698431365
transform -1 0 8400 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _652_
timestamp 1698431365
transform -1 0 15456 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _653_
timestamp 1698431365
transform -1 0 10304 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _654_
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _655_
timestamp 1698431365
transform 1 0 6496 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _656_
timestamp 1698431365
transform 1 0 26320 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _657_
timestamp 1698431365
transform -1 0 8960 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _658_
timestamp 1698431365
transform 1 0 5936 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _659_
timestamp 1698431365
transform 1 0 6496 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _660_
timestamp 1698431365
transform -1 0 9520 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _661_
timestamp 1698431365
transform -1 0 8064 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _662_
timestamp 1698431365
transform 1 0 6608 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _663_
timestamp 1698431365
transform -1 0 27104 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _664_
timestamp 1698431365
transform -1 0 10640 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _665_
timestamp 1698431365
transform 1 0 9184 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _666_
timestamp 1698431365
transform -1 0 10976 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _667_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _668_
timestamp 1698431365
transform -1 0 14000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _669_
timestamp 1698431365
transform -1 0 12768 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _670_
timestamp 1698431365
transform -1 0 12992 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _671_
timestamp 1698431365
transform -1 0 12432 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _672_
timestamp 1698431365
transform -1 0 12096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _673_
timestamp 1698431365
transform 1 0 31808 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _674_
timestamp 1698431365
transform -1 0 14560 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _675_
timestamp 1698431365
transform -1 0 14784 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _676_
timestamp 1698431365
transform -1 0 14112 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _677_
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _678_
timestamp 1698431365
transform 1 0 12544 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _679_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _680_
timestamp 1698431365
transform 1 0 14560 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _681_
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _682_
timestamp 1698431365
transform 1 0 15792 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _683_
timestamp 1698431365
transform 1 0 14560 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _684_
timestamp 1698431365
transform -1 0 18816 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _685_
timestamp 1698431365
transform 1 0 18480 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _686_
timestamp 1698431365
transform -1 0 19040 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _687_
timestamp 1698431365
transform -1 0 21840 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _688_
timestamp 1698431365
transform -1 0 21056 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _689_
timestamp 1698431365
transform 1 0 21392 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _690_
timestamp 1698431365
transform -1 0 19712 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _691_
timestamp 1698431365
transform -1 0 19488 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _692_
timestamp 1698431365
transform -1 0 20384 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _693_
timestamp 1698431365
transform -1 0 20496 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _694_
timestamp 1698431365
transform -1 0 19936 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _695_
timestamp 1698431365
transform -1 0 21392 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _696_
timestamp 1698431365
transform 1 0 20384 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _697_
timestamp 1698431365
transform 1 0 19600 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _698_
timestamp 1698431365
transform -1 0 20832 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _699_
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _700_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _701_
timestamp 1698431365
transform 1 0 21504 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _702_
timestamp 1698431365
transform 1 0 21728 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _703_
timestamp 1698431365
transform 1 0 21840 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _704_
timestamp 1698431365
transform 1 0 19712 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _705_
timestamp 1698431365
transform 1 0 20944 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _706_
timestamp 1698431365
transform -1 0 21616 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _707_
timestamp 1698431365
transform 1 0 19600 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _708_
timestamp 1698431365
transform 1 0 16352 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _709_
timestamp 1698431365
transform -1 0 21056 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _710_
timestamp 1698431365
transform -1 0 18368 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _711_
timestamp 1698431365
transform -1 0 19712 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _712_
timestamp 1698431365
transform 1 0 19152 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _713_
timestamp 1698431365
transform 1 0 18928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _714_
timestamp 1698431365
transform -1 0 20944 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _715_
timestamp 1698431365
transform -1 0 18928 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _716_
timestamp 1698431365
transform 1 0 18368 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _717_
timestamp 1698431365
transform -1 0 20608 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _718_
timestamp 1698431365
transform -1 0 18256 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _719_
timestamp 1698431365
transform 1 0 18144 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _720_
timestamp 1698431365
transform -1 0 18368 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _721_
timestamp 1698431365
transform -1 0 18704 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _722_
timestamp 1698431365
transform -1 0 18144 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _723_
timestamp 1698431365
transform 1 0 22960 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _724_
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _725_
timestamp 1698431365
transform -1 0 29680 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _726_
timestamp 1698431365
transform -1 0 28896 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _727_
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _728_
timestamp 1698431365
transform 1 0 22400 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _729_
timestamp 1698431365
transform 1 0 22064 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _730_
timestamp 1698431365
transform 1 0 23184 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _731_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _732_
timestamp 1698431365
transform 1 0 27328 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _733_
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _734_
timestamp 1698431365
transform 1 0 27888 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _735_
timestamp 1698431365
transform -1 0 28336 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _736_
timestamp 1698431365
transform 1 0 26768 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _737_
timestamp 1698431365
transform 1 0 27104 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _738_
timestamp 1698431365
transform 1 0 27888 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _739_
timestamp 1698431365
transform 1 0 26320 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _740_
timestamp 1698431365
transform 1 0 26768 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _741_
timestamp 1698431365
transform -1 0 29680 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _742_
timestamp 1698431365
transform 1 0 27328 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _743_
timestamp 1698431365
transform 1 0 22288 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _744_
timestamp 1698431365
transform 1 0 23072 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _745_
timestamp 1698431365
transform 1 0 23296 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _746_
timestamp 1698431365
transform 1 0 24864 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _747_
timestamp 1698431365
transform -1 0 27776 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _748_
timestamp 1698431365
transform -1 0 29120 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _749_
timestamp 1698431365
transform 1 0 23520 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _750_
timestamp 1698431365
transform 1 0 26432 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _751_
timestamp 1698431365
transform 1 0 27104 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _752_
timestamp 1698431365
transform 1 0 27664 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _753_
timestamp 1698431365
transform -1 0 27328 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _754_
timestamp 1698431365
transform 1 0 27328 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _755_
timestamp 1698431365
transform 1 0 28000 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _756_
timestamp 1698431365
transform -1 0 25536 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _757_
timestamp 1698431365
transform -1 0 25424 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _758_
timestamp 1698431365
transform -1 0 26656 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _759_
timestamp 1698431365
transform 1 0 27216 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _760_
timestamp 1698431365
transform 1 0 27776 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _761_
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _762_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _763_
timestamp 1698431365
transform 1 0 28896 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _764_
timestamp 1698431365
transform 1 0 33040 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _765_
timestamp 1698431365
transform 1 0 34720 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _766_
timestamp 1698431365
transform 1 0 35168 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _767_
timestamp 1698431365
transform 1 0 33936 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _768_
timestamp 1698431365
transform 1 0 34608 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _769_
timestamp 1698431365
transform 1 0 35280 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _770_
timestamp 1698431365
transform -1 0 36736 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _771_
timestamp 1698431365
transform 1 0 35168 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _772_
timestamp 1698431365
transform -1 0 36624 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _773_
timestamp 1698431365
transform 1 0 34720 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _774_
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _775_
timestamp 1698431365
transform 1 0 29232 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _776_
timestamp 1698431365
transform -1 0 36064 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _777_
timestamp 1698431365
transform 1 0 24528 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _778_
timestamp 1698431365
transform -1 0 24752 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _779_
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _780_
timestamp 1698431365
transform -1 0 23632 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _781_
timestamp 1698431365
transform 1 0 21616 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _782_
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _783_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _784_
timestamp 1698431365
transform -1 0 27776 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _785_
timestamp 1698431365
transform 1 0 26208 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _786_
timestamp 1698431365
transform 1 0 26768 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _787_
timestamp 1698431365
transform 1 0 23856 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _788_
timestamp 1698431365
transform 1 0 22736 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _789_
timestamp 1698431365
transform -1 0 28224 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _790_
timestamp 1698431365
transform 1 0 25872 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _791_
timestamp 1698431365
transform -1 0 28000 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _792_
timestamp 1698431365
transform 1 0 27328 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _793_
timestamp 1698431365
transform 1 0 29120 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _794_
timestamp 1698431365
transform -1 0 30240 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _795_
timestamp 1698431365
transform -1 0 30016 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _796_
timestamp 1698431365
transform 1 0 30016 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _797_
timestamp 1698431365
transform 1 0 29568 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _798_
timestamp 1698431365
transform -1 0 32368 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _799_
timestamp 1698431365
transform 1 0 30128 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _800_
timestamp 1698431365
transform 1 0 30464 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _801_
timestamp 1698431365
transform 1 0 30240 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _802_
timestamp 1698431365
transform 1 0 31024 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _803_
timestamp 1698431365
transform 1 0 23856 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _804_
timestamp 1698431365
transform 1 0 22736 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _805_
timestamp 1698431365
transform 1 0 25088 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _806_
timestamp 1698431365
transform 1 0 29344 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _807_
timestamp 1698431365
transform 1 0 29904 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _808_
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _809_
timestamp 1698431365
transform 1 0 25200 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _810_
timestamp 1698431365
transform -1 0 32256 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _811_
timestamp 1698431365
transform 1 0 30688 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _812_
timestamp 1698431365
transform 1 0 30464 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _813_
timestamp 1698431365
transform 1 0 31248 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _814_
timestamp 1698431365
transform -1 0 31024 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _815_
timestamp 1698431365
transform -1 0 29904 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _816_
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _817_
timestamp 1698431365
transform 1 0 27328 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _818_
timestamp 1698431365
transform -1 0 30128 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _819_
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _820_
timestamp 1698431365
transform 1 0 34048 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _821_
timestamp 1698431365
transform -1 0 36288 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _822_
timestamp 1698431365
transform 1 0 35280 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _823_
timestamp 1698431365
transform -1 0 36064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _824_
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _825_
timestamp 1698431365
transform 1 0 35840 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _826_
timestamp 1698431365
transform 1 0 36064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _827_
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _828_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _829_
timestamp 1698431365
transform 1 0 36176 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _830_
timestamp 1698431365
transform 1 0 35280 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _831_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _832_
timestamp 1698431365
transform -1 0 37744 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _833_
timestamp 1698431365
transform 1 0 32032 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _834_
timestamp 1698431365
transform 1 0 32032 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _835_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38864 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _836_
timestamp 1698431365
transform -1 0 5376 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _837_
timestamp 1698431365
transform -1 0 5152 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _838_
timestamp 1698431365
transform -1 0 5936 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _839_
timestamp 1698431365
transform -1 0 5264 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _840_
timestamp 1698431365
transform -1 0 6048 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _841_
timestamp 1698431365
transform -1 0 5264 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _842_
timestamp 1698431365
transform -1 0 7056 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _843_
timestamp 1698431365
transform -1 0 5040 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _844_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _845_
timestamp 1698431365
transform 1 0 37072 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _846_
timestamp 1698431365
transform 1 0 40320 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _847_
timestamp 1698431365
transform -1 0 8288 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _848_
timestamp 1698431365
transform 1 0 2128 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _849_
timestamp 1698431365
transform 1 0 3584 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _850_
timestamp 1698431365
transform 1 0 1792 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _851_
timestamp 1698431365
transform 1 0 9632 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _852_
timestamp 1698431365
transform -1 0 5040 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _853_
timestamp 1698431365
transform 1 0 11200 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _854_
timestamp 1698431365
transform 1 0 5824 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _855_
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _856_
timestamp 1698431365
transform 1 0 2016 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _857_
timestamp 1698431365
transform 1 0 3136 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _858_
timestamp 1698431365
transform -1 0 9184 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _859_
timestamp 1698431365
transform 1 0 8512 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _860_
timestamp 1698431365
transform 1 0 12432 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _861_
timestamp 1698431365
transform -1 0 14672 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _862_
timestamp 1698431365
transform 1 0 13776 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _863_
timestamp 1698431365
transform 1 0 17136 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _864_
timestamp 1698431365
transform -1 0 20496 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _865_
timestamp 1698431365
transform 1 0 19936 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _866_
timestamp 1698431365
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _867_
timestamp 1698431365
transform 1 0 22736 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _868_
timestamp 1698431365
transform 1 0 23296 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _869_
timestamp 1698431365
transform 1 0 21616 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _870_
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _871_
timestamp 1698431365
transform -1 0 19488 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _872_
timestamp 1698431365
transform -1 0 18144 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _873_
timestamp 1698431365
transform 1 0 21168 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _874_
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _875_
timestamp 1698431365
transform 1 0 27664 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _876_
timestamp 1698431365
transform 1 0 29232 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _877_
timestamp 1698431365
transform 1 0 32480 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _878_
timestamp 1698431365
transform -1 0 24864 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _879_
timestamp 1698431365
transform 1 0 27440 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _880_
timestamp 1698431365
transform 1 0 30912 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _881_
timestamp 1698431365
transform -1 0 28336 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _882_
timestamp 1698431365
transform -1 0 30576 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _883_
timestamp 1698431365
transform 1 0 36288 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _884_
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _885_
timestamp 1698431365
transform 1 0 37296 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _886_
timestamp 1698431365
transform 1 0 38752 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _887_
timestamp 1698431365
transform -1 0 24304 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _888_
timestamp 1698431365
transform -1 0 28896 0 -1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _889_
timestamp 1698431365
transform -1 0 24752 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _890_
timestamp 1698431365
transform -1 0 29456 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _891_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _892_
timestamp 1698431365
transform 1 0 30800 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _893_
timestamp 1698431365
transform 1 0 31808 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _894_
timestamp 1698431365
transform -1 0 24752 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _895_
timestamp 1698431365
transform -1 0 32592 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _896_
timestamp 1698431365
transform 1 0 31808 0 1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _897_
timestamp 1698431365
transform -1 0 34048 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _898_
timestamp 1698431365
transform -1 0 30688 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _899_
timestamp 1698431365
transform 1 0 36176 0 -1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _900_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _901_
timestamp 1698431365
transform 1 0 37072 0 -1 20384
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _902_
timestamp 1698431365
transform 1 0 38080 0 1 20384
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _903_
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _904_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__A1 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__I1
timestamp 1698431365
transform 1 0 17472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__S
timestamp 1698431365
transform 1 0 20496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__I
timestamp 1698431365
transform 1 0 22400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A1
timestamp 1698431365
transform 1 0 23408 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A2
timestamp 1698431365
transform 1 0 24752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__I0
timestamp 1698431365
transform 1 0 29344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__I1
timestamp 1698431365
transform -1 0 30016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__S
timestamp 1698431365
transform 1 0 27216 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__I0
timestamp 1698431365
transform 1 0 32032 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__I1
timestamp 1698431365
transform -1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__S
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__I0
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__I1
timestamp 1698431365
transform -1 0 35504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__S
timestamp 1698431365
transform 1 0 34832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__I0
timestamp 1698431365
transform 1 0 35616 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__I1
timestamp 1698431365
transform -1 0 36736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__S
timestamp 1698431365
transform 1 0 36064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__I
timestamp 1698431365
transform 1 0 22624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A1
timestamp 1698431365
transform 1 0 7168 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A1
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A2
timestamp 1698431365
transform 1 0 14896 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A1
timestamp 1698431365
transform -1 0 12432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A2
timestamp 1698431365
transform -1 0 11536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__A1
timestamp 1698431365
transform -1 0 15456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__A2
timestamp 1698431365
transform 1 0 15680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A1
timestamp 1698431365
transform -1 0 16576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A2
timestamp 1698431365
transform 1 0 14784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__A1
timestamp 1698431365
transform 1 0 8288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__A2
timestamp 1698431365
transform 1 0 7840 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__S
timestamp 1698431365
transform 1 0 37520 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A1
timestamp 1698431365
transform 1 0 30128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A2
timestamp 1698431365
transform 1 0 27440 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__I
timestamp 1698431365
transform 1 0 29680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__A2
timestamp 1698431365
transform -1 0 29904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__I0
timestamp 1698431365
transform 1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__S
timestamp 1698431365
transform 1 0 41104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__I0
timestamp 1698431365
transform 1 0 42112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__S
timestamp 1698431365
transform -1 0 40208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__I0
timestamp 1698431365
transform -1 0 39872 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__S
timestamp 1698431365
transform -1 0 40320 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__I0
timestamp 1698431365
transform 1 0 41216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__S
timestamp 1698431365
transform 1 0 41664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__A1
timestamp 1698431365
transform 1 0 21840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__A2
timestamp 1698431365
transform -1 0 20496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A1
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A1
timestamp 1698431365
transform 1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A2
timestamp 1698431365
transform 1 0 27216 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A1
timestamp 1698431365
transform 1 0 30464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A2
timestamp 1698431365
transform 1 0 29120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__A1
timestamp 1698431365
transform -1 0 32928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__A2
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A1
timestamp 1698431365
transform -1 0 6944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A2
timestamp 1698431365
transform -1 0 6384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A1
timestamp 1698431365
transform -1 0 8624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A2
timestamp 1698431365
transform 1 0 8064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__A2
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A1
timestamp 1698431365
transform -1 0 24304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A2
timestamp 1698431365
transform -1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A2
timestamp 1698431365
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A1
timestamp 1698431365
transform 1 0 29232 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A2
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A1
timestamp 1698431365
transform 1 0 19936 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__I
timestamp 1698431365
transform 1 0 44576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__I
timestamp 1698431365
transform 1 0 11536 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__I
timestamp 1698431365
transform 1 0 35952 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__A1
timestamp 1698431365
transform -1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__A2
timestamp 1698431365
transform -1 0 15232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A2
timestamp 1698431365
transform 1 0 38752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__467__I
timestamp 1698431365
transform -1 0 20608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__I
timestamp 1698431365
transform 1 0 13552 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__I
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__I
timestamp 1698431365
transform 1 0 9744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__I
timestamp 1698431365
transform 1 0 8848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__A3
timestamp 1698431365
transform 1 0 11536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__I
timestamp 1698431365
transform 1 0 17584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__I
timestamp 1698431365
transform -1 0 8064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__I
timestamp 1698431365
transform 1 0 11088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__I
timestamp 1698431365
transform 1 0 10640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__I
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__B2
timestamp 1698431365
transform 1 0 22288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__C2
timestamp 1698431365
transform -1 0 19488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__A1
timestamp 1698431365
transform 1 0 9744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__I
timestamp 1698431365
transform 1 0 18928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A1
timestamp 1698431365
transform 1 0 20384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A2
timestamp 1698431365
transform 1 0 18480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__I
timestamp 1698431365
transform 1 0 7616 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__I
timestamp 1698431365
transform 1 0 8064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__I
timestamp 1698431365
transform -1 0 17920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__I
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A1
timestamp 1698431365
transform 1 0 14896 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A2
timestamp 1698431365
transform 1 0 16016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__B2
timestamp 1698431365
transform 1 0 13216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__C
timestamp 1698431365
transform 1 0 8512 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A1
timestamp 1698431365
transform -1 0 9856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A2
timestamp 1698431365
transform 1 0 9856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__A2
timestamp 1698431365
transform 1 0 15680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__C1
timestamp 1698431365
transform -1 0 16352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__I
timestamp 1698431365
transform 1 0 17808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__I
timestamp 1698431365
transform 1 0 17584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A1
timestamp 1698431365
transform -1 0 20384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__C
timestamp 1698431365
transform -1 0 8400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A1
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__B2
timestamp 1698431365
transform 1 0 17584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__I
timestamp 1698431365
transform 1 0 15680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__I
timestamp 1698431365
transform 1 0 13216 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__A1
timestamp 1698431365
transform 1 0 12432 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__C1
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__I
timestamp 1698431365
transform 1 0 18032 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A1
timestamp 1698431365
transform -1 0 11536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A2
timestamp 1698431365
transform 1 0 10752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__B2
timestamp 1698431365
transform -1 0 8400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__I
timestamp 1698431365
transform 1 0 15456 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__A1
timestamp 1698431365
transform 1 0 19936 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__B2
timestamp 1698431365
transform 1 0 20384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__C2
timestamp 1698431365
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__A2
timestamp 1698431365
transform 1 0 14672 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__B1
timestamp 1698431365
transform 1 0 19824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__B2
timestamp 1698431365
transform -1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__C1
timestamp 1698431365
transform 1 0 20272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A1
timestamp 1698431365
transform 1 0 13104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__A1
timestamp 1698431365
transform -1 0 17248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__B2
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__554__A1
timestamp 1698431365
transform -1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__554__B2
timestamp 1698431365
transform -1 0 14336 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__B1
timestamp 1698431365
transform -1 0 13664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__B2
timestamp 1698431365
transform -1 0 13776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__C1
timestamp 1698431365
transform 1 0 13888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__A1
timestamp 1698431365
transform 1 0 19712 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__A1
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__B2
timestamp 1698431365
transform -1 0 17920 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__C2
timestamp 1698431365
transform -1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__A1
timestamp 1698431365
transform -1 0 12992 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__A1
timestamp 1698431365
transform -1 0 14112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__A2
timestamp 1698431365
transform 1 0 14784 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__B2
timestamp 1698431365
transform 1 0 14336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__563__A1
timestamp 1698431365
transform 1 0 11088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__A1
timestamp 1698431365
transform 1 0 18480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__B2
timestamp 1698431365
transform 1 0 17024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__A1
timestamp 1698431365
transform -1 0 17472 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__B2
timestamp 1698431365
transform 1 0 15904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__C2
timestamp 1698431365
transform -1 0 14112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__569__B2
timestamp 1698431365
transform 1 0 16800 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__569__C1
timestamp 1698431365
transform -1 0 17472 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__570__A1
timestamp 1698431365
transform 1 0 19936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__571__A1
timestamp 1698431365
transform -1 0 19152 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__571__B2
timestamp 1698431365
transform -1 0 20608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__C
timestamp 1698431365
transform 1 0 10864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__577__C
timestamp 1698431365
transform 1 0 14560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__A1
timestamp 1698431365
transform 1 0 18032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__B2
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__579__B2
timestamp 1698431365
transform 1 0 10416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A1
timestamp 1698431365
transform -1 0 16576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__A1
timestamp 1698431365
transform 1 0 22736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__B2
timestamp 1698431365
transform 1 0 23184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__C1
timestamp 1698431365
transform 1 0 19488 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__583__C
timestamp 1698431365
transform 1 0 10192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__I
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A1
timestamp 1698431365
transform 1 0 21952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A2
timestamp 1698431365
transform 1 0 23296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__A1
timestamp 1698431365
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__A3
timestamp 1698431365
transform 1 0 32816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__A2
timestamp 1698431365
transform 1 0 22848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__A1
timestamp 1698431365
transform 1 0 35728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__593__I
timestamp 1698431365
transform 1 0 29792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__A1
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__A3
timestamp 1698431365
transform -1 0 33824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__A2
timestamp 1698431365
transform -1 0 31360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__597__A1
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__I
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A1
timestamp 1698431365
transform 1 0 34048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A3
timestamp 1698431365
transform 1 0 34048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__601__A2
timestamp 1698431365
transform 1 0 39536 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A1
timestamp 1698431365
transform -1 0 40208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__I
timestamp 1698431365
transform 1 0 16128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__A1
timestamp 1698431365
transform 1 0 19376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__A2
timestamp 1698431365
transform 1 0 20384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__609__A1
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__611__A2
timestamp 1698431365
transform -1 0 10528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__615__I
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__A1
timestamp 1698431365
transform -1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__620__C
timestamp 1698431365
transform 1 0 4480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__621__I
timestamp 1698431365
transform 1 0 23744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__622__A1
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__A1
timestamp 1698431365
transform 1 0 3360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__C
timestamp 1698431365
transform -1 0 4928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__I
timestamp 1698431365
transform 1 0 25648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__630__A1
timestamp 1698431365
transform -1 0 11648 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__A1
timestamp 1698431365
transform 1 0 4928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__635__I
timestamp 1698431365
transform 1 0 35168 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__637__C
timestamp 1698431365
transform 1 0 6832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__I
timestamp 1698431365
transform 1 0 25312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__639__A1
timestamp 1698431365
transform -1 0 13776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__642__I
timestamp 1698431365
transform 1 0 20384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__643__A1
timestamp 1698431365
transform 1 0 14336 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__645__I
timestamp 1698431365
transform 1 0 11424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__B
timestamp 1698431365
transform -1 0 9408 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__649__A2
timestamp 1698431365
transform -1 0 16800 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__A1
timestamp 1698431365
transform 1 0 8624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__A2
timestamp 1698431365
transform -1 0 16352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__654__A1
timestamp 1698431365
transform -1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__B
timestamp 1698431365
transform 1 0 7728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__I
timestamp 1698431365
transform 1 0 26096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__A1
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__B
timestamp 1698431365
transform 1 0 7616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__660__A1
timestamp 1698431365
transform 1 0 9744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__661__A1
timestamp 1698431365
transform -1 0 7504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__662__B
timestamp 1698431365
transform 1 0 7616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__663__I
timestamp 1698431365
transform 1 0 25984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__664__A1
timestamp 1698431365
transform 1 0 10864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__665__A1
timestamp 1698431365
transform 1 0 8960 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__669__A1
timestamp 1698431365
transform 1 0 11984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__671__A1
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__I
timestamp 1698431365
transform -1 0 31808 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__A1
timestamp 1698431365
transform -1 0 14000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__A1
timestamp 1698431365
transform 1 0 14784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__A1
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__A1
timestamp 1698431365
transform -1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__A1
timestamp 1698431365
transform 1 0 14336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__A1
timestamp 1698431365
transform 1 0 18256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__A1
timestamp 1698431365
transform -1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__690__A1
timestamp 1698431365
transform -1 0 20160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__692__I
timestamp 1698431365
transform 1 0 18592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__693__A1
timestamp 1698431365
transform 1 0 19600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__694__C
timestamp 1698431365
transform -1 0 20160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__A1
timestamp 1698431365
transform -1 0 20720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__696__A1
timestamp 1698431365
transform 1 0 22176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__696__C
timestamp 1698431365
transform 1 0 21728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__697__A1
timestamp 1698431365
transform 1 0 19376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__699__A1
timestamp 1698431365
transform 1 0 20832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__A1
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__702__A1
timestamp 1698431365
transform 1 0 23520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__702__C
timestamp 1698431365
transform 1 0 23072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__703__A1
timestamp 1698431365
transform 1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__704__A1
timestamp 1698431365
transform -1 0 19712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__706__A1
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__A1
timestamp 1698431365
transform 1 0 19376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__B
timestamp 1698431365
transform -1 0 20160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__A1
timestamp 1698431365
transform 1 0 17584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__A1
timestamp 1698431365
transform 1 0 19936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__B
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__A1
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__A2
timestamp 1698431365
transform 1 0 20048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__A1
timestamp 1698431365
transform -1 0 17808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__A2
timestamp 1698431365
transform 1 0 19152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__B
timestamp 1698431365
transform -1 0 19488 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__A1
timestamp 1698431365
transform -1 0 19376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__B
timestamp 1698431365
transform -1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__A1
timestamp 1698431365
transform 1 0 23744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__A1
timestamp 1698431365
transform 1 0 21392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__725__I
timestamp 1698431365
transform 1 0 29904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__728__A1
timestamp 1698431365
transform -1 0 22400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__A1
timestamp 1698431365
transform 1 0 22848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__A1
timestamp 1698431365
transform 1 0 26544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__A1
timestamp 1698431365
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__736__A1
timestamp 1698431365
transform 1 0 26544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__A1
timestamp 1698431365
transform -1 0 28896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__739__A1
timestamp 1698431365
transform 1 0 26096 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__A1
timestamp 1698431365
transform 1 0 29120 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__743__A1
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__746__A1
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__746__A2
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__748__A1
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__749__A1
timestamp 1698431365
transform 1 0 23296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__753__A1
timestamp 1698431365
transform 1 0 26544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__756__A1
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__758__A1
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__759__A1
timestamp 1698431365
transform 1 0 26992 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__760__A1
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__763__A1
timestamp 1698431365
transform 1 0 29680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__765__A1
timestamp 1698431365
transform 1 0 34496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__767__A1
timestamp 1698431365
transform 1 0 33712 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__768__A1
timestamp 1698431365
transform 1 0 34384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__770__A1
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__771__A1
timestamp 1698431365
transform 1 0 36848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__773__A1
timestamp 1698431365
transform 1 0 34496 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__774__A1
timestamp 1698431365
transform 1 0 37968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__776__B
timestamp 1698431365
transform -1 0 35168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__777__A1
timestamp 1698431365
transform 1 0 25312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__780__A1
timestamp 1698431365
transform 1 0 22736 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__781__A1
timestamp 1698431365
transform 1 0 22288 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__782__A1
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__782__A2
timestamp 1698431365
transform 1 0 24192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__784__A1
timestamp 1698431365
transform 1 0 26992 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__785__A1
timestamp 1698431365
transform 1 0 26992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__786__B
timestamp 1698431365
transform 1 0 27888 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__787__A1
timestamp 1698431365
transform 1 0 22512 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__788__A1
timestamp 1698431365
transform 1 0 25312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__789__A1
timestamp 1698431365
transform 1 0 28448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__791__A1
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__792__B
timestamp 1698431365
transform -1 0 28672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__793__A1
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__794__A1
timestamp 1698431365
transform 1 0 31024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__795__B
timestamp 1698431365
transform -1 0 30464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__796__A1
timestamp 1698431365
transform -1 0 30016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__797__A1
timestamp 1698431365
transform 1 0 29344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__800__A1
timestamp 1698431365
transform -1 0 30464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__801__A1
timestamp 1698431365
transform 1 0 31472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__803__A1
timestamp 1698431365
transform 1 0 23856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__805__A1
timestamp 1698431365
transform 1 0 25872 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__805__A2
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__807__A1
timestamp 1698431365
transform 1 0 29680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__808__C
timestamp 1698431365
transform 1 0 31472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__809__A1
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__809__A2
timestamp 1698431365
transform 1 0 24528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__811__A1
timestamp 1698431365
transform 1 0 31472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__812__A1
timestamp 1698431365
transform 1 0 31248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__814__A1
timestamp 1698431365
transform 1 0 30240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__815__A1
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__817__A1
timestamp 1698431365
transform 1 0 27104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__818__C
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__819__A1
timestamp 1698431365
transform -1 0 31248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__821__A1
timestamp 1698431365
transform 1 0 37184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__824__A1
timestamp 1698431365
transform 1 0 33712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__825__A1
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__827__A1
timestamp 1698431365
transform 1 0 34496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__828__A1
timestamp 1698431365
transform 1 0 35840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__830__A1
timestamp 1698431365
transform -1 0 35280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__831__A1
timestamp 1698431365
transform 1 0 38080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__833__A1
timestamp 1698431365
transform 1 0 31808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__834__A1
timestamp 1698431365
transform -1 0 32032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__835__CLK
timestamp 1698431365
transform 1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__836__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__837__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__838__CLK
timestamp 1698431365
transform -1 0 6384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__839__CLK
timestamp 1698431365
transform -1 0 5936 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__840__CLK
timestamp 1698431365
transform 1 0 6272 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__841__CLK
timestamp 1698431365
transform 1 0 5712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__842__CLK
timestamp 1698431365
transform 1 0 7280 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__843__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__844__CLK
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__845__CLK
timestamp 1698431365
transform 1 0 36176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__846__CLK
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__847__CLK
timestamp 1698431365
transform 1 0 8512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__848__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__849__CLK
timestamp 1698431365
transform 1 0 6832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__850__CLK
timestamp 1698431365
transform 1 0 5712 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__851__CLK
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__852__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__853__CLK
timestamp 1698431365
transform -1 0 14896 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__854__CLK
timestamp 1698431365
transform 1 0 9296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__855__CLK
timestamp 1698431365
transform -1 0 5936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__856__CLK
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__857__CLK
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__858__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__859__CLK
timestamp 1698431365
transform 1 0 11760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__860__CLK
timestamp 1698431365
transform 1 0 15904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__861__CLK
timestamp 1698431365
transform 1 0 14784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__862__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__863__CLK
timestamp 1698431365
transform 1 0 16912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__864__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__865__CLK
timestamp 1698431365
transform 1 0 19712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__866__CLK
timestamp 1698431365
transform -1 0 21616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__867__CLK
timestamp 1698431365
transform -1 0 26432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__868__CLK
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__869__CLK
timestamp 1698431365
transform -1 0 25536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__870__CLK
timestamp 1698431365
transform 1 0 18144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__871__CLK
timestamp 1698431365
transform 1 0 19712 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__872__CLK
timestamp 1698431365
transform 1 0 18480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__873__CLK
timestamp 1698431365
transform 1 0 21840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__874__CLK
timestamp 1698431365
transform -1 0 28784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__875__CLK
timestamp 1698431365
transform 1 0 31136 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__876__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__877__CLK
timestamp 1698431365
transform 1 0 35952 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__878__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__879__CLK
timestamp 1698431365
transform 1 0 30912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__880__CLK
timestamp 1698431365
transform 1 0 34384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__881__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__882__CLK
timestamp 1698431365
transform -1 0 31024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__883__CLK
timestamp 1698431365
transform 1 0 36064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__884__CLK
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__885__CLK
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__886__CLK
timestamp 1698431365
transform 1 0 38528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__887__CLK
timestamp 1698431365
transform 1 0 24528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__888__CLK
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__889__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__890__CLK
timestamp 1698431365
transform 1 0 29680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__891__CLK
timestamp 1698431365
transform 1 0 32704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__892__CLK
timestamp 1698431365
transform 1 0 34496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__893__CLK
timestamp 1698431365
transform 1 0 31584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__894__CLK
timestamp 1698431365
transform 1 0 25984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__895__CLK
timestamp 1698431365
transform -1 0 33376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__896__CLK
timestamp 1698431365
transform 1 0 35504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__897__CLK
timestamp 1698431365
transform 1 0 34944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__898__CLK
timestamp 1698431365
transform -1 0 31136 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__899__CLK
timestamp 1698431365
transform 1 0 39872 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__900__CLK
timestamp 1698431365
transform 1 0 37632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__901__CLK
timestamp 1698431365
transform 1 0 37632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__902__CLK
timestamp 1698431365
transform 1 0 37856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__903__CLK
timestamp 1698431365
transform 1 0 32704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__904__CLK
timestamp 1698431365
transform 1 0 37072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 27216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 21616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 28896 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 32704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 20272 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 30800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 47712 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 47712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 47712 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 47712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 2912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 2464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 1792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 37072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 1792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 1792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 1792 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 1792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 1792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 6608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 16352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 17696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 18928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 20160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 21616 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 22960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 4704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 5376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 7168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 8176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 9632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 10864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 12768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 13552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 14896 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 47712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 47712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 47712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 47040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 47712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 47712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1698431365
transform 1 0 28448 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output64_I
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output65_I
timestamp 1698431365
transform 1 0 22064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output83_I
timestamp 1698431365
transform 1 0 42784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output84_I
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output85_I
timestamp 1698431365
transform 1 0 46592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1698431365
transform -1 0 20048 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1698431365
transform 1 0 31024 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_40 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_74
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_108
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_165
timestamp 1698431365
transform 1 0 19824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_300
timestamp 1698431365
transform 1 0 34944 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_314
timestamp 1698431365
transform 1 0 36512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_316
timestamp 1698431365
transform 1 0 36736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_325 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37744 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_333
timestamp 1698431365
transform 1 0 38640 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_337
timestamp 1698431365
transform 1 0 39088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_368
timestamp 1698431365
transform 1 0 42560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_372
timestamp 1698431365
transform 1 0 43008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_402
timestamp 1698431365
transform 1 0 46368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_406
timestamp 1698431365
transform 1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698431365
transform 1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_8
timestamp 1698431365
transform 1 0 2240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_12
timestamp 1698431365
transform 1 0 2688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_16
timestamp 1698431365
transform 1 0 3136 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_24
timestamp 1698431365
transform 1 0 4032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_28
timestamp 1698431365
transform 1 0 4480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_30
timestamp 1698431365
transform 1 0 4704 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_57
timestamp 1698431365
transform 1 0 7728 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_65
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_98
timestamp 1698431365
transform 1 0 12320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_102
timestamp 1698431365
transform 1 0 12768 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_129
timestamp 1698431365
transform 1 0 15792 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_137
timestamp 1698431365
transform 1 0 16688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698431365
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_183
timestamp 1698431365
transform 1 0 21840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_187 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_228
timestamp 1698431365
transform 1 0 26880 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_255
timestamp 1698431365
transform 1 0 29904 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_271
timestamp 1698431365
transform 1 0 31696 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_309 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35952 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_341
timestamp 1698431365
transform 1 0 39536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_345
timestamp 1698431365
transform 1 0 39984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_347
timestamp 1698431365
transform 1 0 40208 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_354
timestamp 1698431365
transform 1 0 40992 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_381
timestamp 1698431365
transform 1 0 44016 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_397
timestamp 1698431365
transform 1 0 45808 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_405
timestamp 1698431365
transform 1 0 46704 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_408
timestamp 1698431365
transform 1 0 47040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_6
timestamp 1698431365
transform 1 0 2016 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698431365
transform 1 0 3808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698431365
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_185
timestamp 1698431365
transform 1 0 22064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_219
timestamp 1698431365
transform 1 0 25872 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_235
timestamp 1698431365
transform 1 0 27664 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_419
timestamp 1698431365
transform 1 0 48272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_10
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_42
timestamp 1698431365
transform 1 0 6048 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_58
timestamp 1698431365
transform 1 0 7840 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_158
timestamp 1698431365
transform 1 0 19040 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_162
timestamp 1698431365
transform 1 0 19488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_195
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_207
timestamp 1698431365
transform 1 0 24528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_139
timestamp 1698431365
transform 1 0 16912 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_155
timestamp 1698431365
transform 1 0 18704 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_163
timestamp 1698431365
transform 1 0 19600 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_167
timestamp 1698431365
transform 1 0 20048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_201
timestamp 1698431365
transform 1 0 23856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_205
timestamp 1698431365
transform 1 0 24304 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_237
timestamp 1698431365
transform 1 0 27888 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_419
timestamp 1698431365
transform 1 0 48272 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_8
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_12
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_60
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_181
timestamp 1698431365
transform 1 0 21616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_185
timestamp 1698431365
transform 1 0 22064 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_155
timestamp 1698431365
transform 1 0 18704 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_163
timestamp 1698431365
transform 1 0 19600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_165
timestamp 1698431365
transform 1 0 19824 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_168
timestamp 1698431365
transform 1 0 20160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_185
timestamp 1698431365
transform 1 0 22064 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_220
timestamp 1698431365
transform 1 0 25984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_224
timestamp 1698431365
transform 1 0 26432 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_419
timestamp 1698431365
transform 1 0 48272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_12
timestamp 1698431365
transform 1 0 2688 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_44
timestamp 1698431365
transform 1 0 6272 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_60
timestamp 1698431365
transform 1 0 8064 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_88
timestamp 1698431365
transform 1 0 11200 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_91
timestamp 1698431365
transform 1 0 11536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_95
timestamp 1698431365
transform 1 0 11984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_128
timestamp 1698431365
transform 1 0 15680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_132
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_180
timestamp 1698431365
transform 1 0 21504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_184
timestamp 1698431365
transform 1 0 21952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_188
timestamp 1698431365
transform 1 0 22400 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_204
timestamp 1698431365
transform 1 0 24192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_208
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_216
timestamp 1698431365
transform 1 0 25536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_228
timestamp 1698431365
transform 1 0 26880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_232
timestamp 1698431365
transform 1 0 27328 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_264
timestamp 1698431365
transform 1 0 30912 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_384
timestamp 1698431365
transform 1 0 44352 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_400
timestamp 1698431365
transform 1 0 46144 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_408
timestamp 1698431365
transform 1 0 47040 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_6
timestamp 1698431365
transform 1 0 2016 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_22
timestamp 1698431365
transform 1 0 3808 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_30
timestamp 1698431365
transform 1 0 4704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_63
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698431365
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_118
timestamp 1698431365
transform 1 0 14560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_122
timestamp 1698431365
transform 1 0 15008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_126
timestamp 1698431365
transform 1 0 15456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_130
timestamp 1698431365
transform 1 0 15904 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_162
timestamp 1698431365
transform 1 0 19488 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_192
timestamp 1698431365
transform 1 0 22848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_196
timestamp 1698431365
transform 1 0 23296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_200
timestamp 1698431365
transform 1 0 23744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_208
timestamp 1698431365
transform 1 0 24640 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_240
timestamp 1698431365
transform 1 0 28224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_278
timestamp 1698431365
transform 1 0 32480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_282
timestamp 1698431365
transform 1 0 32928 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_419
timestamp 1698431365
transform 1 0 48272 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_10
timestamp 1698431365
transform 1 0 2464 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_42
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_119
timestamp 1698431365
transform 1 0 14672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_133
timestamp 1698431365
transform 1 0 16240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_164
timestamp 1698431365
transform 1 0 19712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_168
timestamp 1698431365
transform 1 0 20160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_170
timestamp 1698431365
transform 1 0 20384 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_185
timestamp 1698431365
transform 1 0 22064 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_201
timestamp 1698431365
transform 1 0 23856 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_251
timestamp 1698431365
transform 1 0 29456 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_255
timestamp 1698431365
transform 1 0 29904 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_271
timestamp 1698431365
transform 1 0 31696 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_6
timestamp 1698431365
transform 1 0 2016 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_22
timestamp 1698431365
transform 1 0 3808 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_30
timestamp 1698431365
transform 1 0 4704 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_115
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_119
timestamp 1698431365
transform 1 0 14672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_132
timestamp 1698431365
transform 1 0 16128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_136
timestamp 1698431365
transform 1 0 16576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_138
timestamp 1698431365
transform 1 0 16800 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_170
timestamp 1698431365
transform 1 0 20384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_179
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_186
timestamp 1698431365
transform 1 0 22176 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_218
timestamp 1698431365
transform 1 0 25760 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_234
timestamp 1698431365
transform 1 0 27552 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698431365
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_294
timestamp 1698431365
transform 1 0 34272 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_298
timestamp 1698431365
transform 1 0 34720 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_419
timestamp 1698431365
transform 1 0 48272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_26
timestamp 1698431365
transform 1 0 4256 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_38
timestamp 1698431365
transform 1 0 5600 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_76
timestamp 1698431365
transform 1 0 9856 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_99
timestamp 1698431365
transform 1 0 12432 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_103
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_105
timestamp 1698431365
transform 1 0 13104 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_114
timestamp 1698431365
transform 1 0 14112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_118
timestamp 1698431365
transform 1 0 14560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_176
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_228
timestamp 1698431365
transform 1 0 26880 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_240
timestamp 1698431365
transform 1 0 28224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_244
timestamp 1698431365
transform 1 0 28672 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_256
timestamp 1698431365
transform 1 0 30016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_260
timestamp 1698431365
transform 1 0 30464 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_268
timestamp 1698431365
transform 1 0 31360 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_272
timestamp 1698431365
transform 1 0 31808 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_6
timestamp 1698431365
transform 1 0 2016 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_22
timestamp 1698431365
transform 1 0 3808 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_85
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_87
timestamp 1698431365
transform 1 0 11088 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_96
timestamp 1698431365
transform 1 0 12096 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_120
timestamp 1698431365
transform 1 0 14784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_122
timestamp 1698431365
transform 1 0 15008 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_195
timestamp 1698431365
transform 1 0 23184 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_225
timestamp 1698431365
transform 1 0 26544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_229
timestamp 1698431365
transform 1 0 26992 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698431365
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_263
timestamp 1698431365
transform 1 0 30800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_267
timestamp 1698431365
transform 1 0 31248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_271
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_303
timestamp 1698431365
transform 1 0 35280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_419
timestamp 1698431365
transform 1 0 48272 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_10
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_42
timestamp 1698431365
transform 1 0 6048 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_58
timestamp 1698431365
transform 1 0 7840 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_86
timestamp 1698431365
transform 1 0 10976 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_92
timestamp 1698431365
transform 1 0 11648 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_124
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_176
timestamp 1698431365
transform 1 0 21056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_178
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_228
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_230
timestamp 1698431365
transform 1 0 27104 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_233
timestamp 1698431365
transform 1 0 27440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_240
timestamp 1698431365
transform 1 0 28224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_244
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_248
timestamp 1698431365
transform 1 0 29120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_273
timestamp 1698431365
transform 1 0 31920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698431365
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_10
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_41
timestamp 1698431365
transform 1 0 5936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_61
timestamp 1698431365
transform 1 0 8176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_65
timestamp 1698431365
transform 1 0 8624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_67
timestamp 1698431365
transform 1 0 8848 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_75
timestamp 1698431365
transform 1 0 9744 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_83
timestamp 1698431365
transform 1 0 10640 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_90
timestamp 1698431365
transform 1 0 11424 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_94
timestamp 1698431365
transform 1 0 11872 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_102
timestamp 1698431365
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_126
timestamp 1698431365
transform 1 0 15456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_128
timestamp 1698431365
transform 1 0 15680 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_135
timestamp 1698431365
transform 1 0 16464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_158
timestamp 1698431365
transform 1 0 19040 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_297
timestamp 1698431365
transform 1 0 34608 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_313
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_403
timestamp 1698431365
transform 1 0 46480 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_411
timestamp 1698431365
transform 1 0 47376 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_6
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_46
timestamp 1698431365
transform 1 0 6496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_50
timestamp 1698431365
transform 1 0 6944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_52
timestamp 1698431365
transform 1 0 7168 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_55
timestamp 1698431365
transform 1 0 7504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_59
timestamp 1698431365
transform 1 0 7952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_67
timestamp 1698431365
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_83
timestamp 1698431365
transform 1 0 10640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_87
timestamp 1698431365
transform 1 0 11088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_95
timestamp 1698431365
transform 1 0 11984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_97
timestamp 1698431365
transform 1 0 12208 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_109
timestamp 1698431365
transform 1 0 13552 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_146
timestamp 1698431365
transform 1 0 17696 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_154
timestamp 1698431365
transform 1 0 18592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_160
timestamp 1698431365
transform 1 0 19264 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_188
timestamp 1698431365
transform 1 0 22400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_230
timestamp 1698431365
transform 1 0 27104 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_238
timestamp 1698431365
transform 1 0 28000 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_242
timestamp 1698431365
transform 1 0 28448 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_245
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_253
timestamp 1698431365
transform 1 0 29680 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_261
timestamp 1698431365
transform 1 0 30576 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_269
timestamp 1698431365
transform 1 0 31472 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_306
timestamp 1698431365
transform 1 0 35616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_310
timestamp 1698431365
transform 1 0 36064 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_342
timestamp 1698431365
transform 1 0 39648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_6
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_22
timestamp 1698431365
transform 1 0 3808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_30
timestamp 1698431365
transform 1 0 4704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_54
timestamp 1698431365
transform 1 0 7392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_63
timestamp 1698431365
transform 1 0 8400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_67
timestamp 1698431365
transform 1 0 8848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_71
timestamp 1698431365
transform 1 0 9296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_73
timestamp 1698431365
transform 1 0 9520 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_80
timestamp 1698431365
transform 1 0 10304 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_96
timestamp 1698431365
transform 1 0 12096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_100
timestamp 1698431365
transform 1 0 12544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_102
timestamp 1698431365
transform 1 0 12768 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_113
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_128
timestamp 1698431365
transform 1 0 15680 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_150
timestamp 1698431365
transform 1 0 18144 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1698431365
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_183
timestamp 1698431365
transform 1 0 21840 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_215
timestamp 1698431365
transform 1 0 25424 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_231
timestamp 1698431365
transform 1 0 27216 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_239
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_303
timestamp 1698431365
transform 1 0 35280 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_348
timestamp 1698431365
transform 1 0 40320 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_380
timestamp 1698431365
transform 1 0 43904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_419
timestamp 1698431365
transform 1 0 48272 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_45
timestamp 1698431365
transform 1 0 6384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_60
timestamp 1698431365
transform 1 0 8064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_62
timestamp 1698431365
transform 1 0 8288 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_65
timestamp 1698431365
transform 1 0 8624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_67
timestamp 1698431365
transform 1 0 8848 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_80
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_120
timestamp 1698431365
transform 1 0 14784 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_152
timestamp 1698431365
transform 1 0 18368 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_159
timestamp 1698431365
transform 1 0 19152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_250
timestamp 1698431365
transform 1 0 29344 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_260
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_267
timestamp 1698431365
transform 1 0 31248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_271
timestamp 1698431365
transform 1 0 31696 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_287
timestamp 1698431365
transform 1 0 33488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_291
timestamp 1698431365
transform 1 0 33936 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_299
timestamp 1698431365
transform 1 0 34832 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_301
timestamp 1698431365
transform 1 0 35056 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_318
timestamp 1698431365
transform 1 0 36960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_322
timestamp 1698431365
transform 1 0 37408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_326
timestamp 1698431365
transform 1 0 37856 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_342
timestamp 1698431365
transform 1 0 39648 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698431365
transform 1 0 9520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_77
timestamp 1698431365
transform 1 0 9968 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_157
timestamp 1698431365
transform 1 0 18928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_167
timestamp 1698431365
transform 1 0 20048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_209
timestamp 1698431365
transform 1 0 24752 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_213
timestamp 1698431365
transform 1 0 25200 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_224
timestamp 1698431365
transform 1 0 26432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_228
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_238
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_249
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_265
timestamp 1698431365
transform 1 0 31024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_275
timestamp 1698431365
transform 1 0 32144 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_279
timestamp 1698431365
transform 1 0 32592 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_282
timestamp 1698431365
transform 1 0 32928 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_298
timestamp 1698431365
transform 1 0 34720 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_306
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_321
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_419
timestamp 1698431365
transform 1 0 48272 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_12
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_28
timestamp 1698431365
transform 1 0 4480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_36
timestamp 1698431365
transform 1 0 5376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_50
timestamp 1698431365
transform 1 0 6944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_54
timestamp 1698431365
transform 1 0 7392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_58
timestamp 1698431365
transform 1 0 7840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_62
timestamp 1698431365
transform 1 0 8288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_74
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_77
timestamp 1698431365
transform 1 0 9968 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_81
timestamp 1698431365
transform 1 0 10416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_85
timestamp 1698431365
transform 1 0 10864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_89
timestamp 1698431365
transform 1 0 11312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_130
timestamp 1698431365
transform 1 0 15904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1698431365
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_181
timestamp 1698431365
transform 1 0 21616 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_197
timestamp 1698431365
transform 1 0 23408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_199
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_252
timestamp 1698431365
transform 1 0 29568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_256
timestamp 1698431365
transform 1 0 30016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_262
timestamp 1698431365
transform 1 0 30688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_266
timestamp 1698431365
transform 1 0 31136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_332
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_348
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_53
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_65
timestamp 1698431365
transform 1 0 8624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_109
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_118
timestamp 1698431365
transform 1 0 14560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_120
timestamp 1698431365
transform 1 0 14784 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_134
timestamp 1698431365
transform 1 0 16352 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_138
timestamp 1698431365
transform 1 0 16800 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_146
timestamp 1698431365
transform 1 0 17696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_152
timestamp 1698431365
transform 1 0 18368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_156
timestamp 1698431365
transform 1 0 18816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_158
timestamp 1698431365
transform 1 0 19040 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_164
timestamp 1698431365
transform 1 0 19712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_168
timestamp 1698431365
transform 1 0 20160 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_209
timestamp 1698431365
transform 1 0 24752 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_225
timestamp 1698431365
transform 1 0 26544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_235
timestamp 1698431365
transform 1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_239
timestamp 1698431365
transform 1 0 28112 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_259
timestamp 1698431365
transform 1 0 30352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_265
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_269
timestamp 1698431365
transform 1 0 31472 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_276
timestamp 1698431365
transform 1 0 32256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_282
timestamp 1698431365
transform 1 0 32928 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_298
timestamp 1698431365
transform 1 0 34720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_300
timestamp 1698431365
transform 1 0 34944 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_303
timestamp 1698431365
transform 1 0 35280 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_307
timestamp 1698431365
transform 1 0 35728 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_322
timestamp 1698431365
transform 1 0 37408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_326
timestamp 1698431365
transform 1 0 37856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_330
timestamp 1698431365
transform 1 0 38304 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_362
timestamp 1698431365
transform 1 0 41888 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_378
timestamp 1698431365
transform 1 0 43680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_382
timestamp 1698431365
transform 1 0 44128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_419
timestamp 1698431365
transform 1 0 48272 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_44
timestamp 1698431365
transform 1 0 6272 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_52
timestamp 1698431365
transform 1 0 7168 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_56
timestamp 1698431365
transform 1 0 7616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_60
timestamp 1698431365
transform 1 0 8064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_74
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_158
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_166
timestamp 1698431365
transform 1 0 19936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_180
timestamp 1698431365
transform 1 0 21504 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_188
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_194
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_198
timestamp 1698431365
transform 1 0 23520 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_202
timestamp 1698431365
transform 1 0 23968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_227
timestamp 1698431365
transform 1 0 26768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_231
timestamp 1698431365
transform 1 0 27216 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_247
timestamp 1698431365
transform 1 0 29008 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_255
timestamp 1698431365
transform 1 0 29904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_257
timestamp 1698431365
transform 1 0 30128 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_265
timestamp 1698431365
transform 1 0 31024 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_269
timestamp 1698431365
transform 1 0 31472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_290
timestamp 1698431365
transform 1 0 33824 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_294
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_308
timestamp 1698431365
transform 1 0 35840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_310
timestamp 1698431365
transform 1 0 36064 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_384
timestamp 1698431365
transform 1 0 44352 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_400
timestamp 1698431365
transform 1 0 46144 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_408
timestamp 1698431365
transform 1 0 47040 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_87
timestamp 1698431365
transform 1 0 11088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_150
timestamp 1698431365
transform 1 0 18144 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_166
timestamp 1698431365
transform 1 0 19936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_183
timestamp 1698431365
transform 1 0 21840 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_202
timestamp 1698431365
transform 1 0 23968 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_206
timestamp 1698431365
transform 1 0 24416 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_209
timestamp 1698431365
transform 1 0 24752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_221
timestamp 1698431365
transform 1 0 26096 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_237
timestamp 1698431365
transform 1 0 27888 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_249
timestamp 1698431365
transform 1 0 29232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_298
timestamp 1698431365
transform 1 0 34720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_302
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698431365
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_327
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_359
timestamp 1698431365
transform 1 0 41552 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_375
timestamp 1698431365
transform 1 0 43344 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_419
timestamp 1698431365
transform 1 0 48272 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_40
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_58
timestamp 1698431365
transform 1 0 7840 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_158
timestamp 1698431365
transform 1 0 19040 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_160
timestamp 1698431365
transform 1 0 19264 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_168
timestamp 1698431365
transform 1 0 20160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_183
timestamp 1698431365
transform 1 0 21840 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_203
timestamp 1698431365
transform 1 0 24080 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_207
timestamp 1698431365
transform 1 0 24528 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_300
timestamp 1698431365
transform 1 0 34944 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_304
timestamp 1698431365
transform 1 0 35392 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_320
timestamp 1698431365
transform 1 0 37184 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_324
timestamp 1698431365
transform 1 0 37632 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_328
timestamp 1698431365
transform 1 0 38080 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_344
timestamp 1698431365
transform 1 0 39872 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_348
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_4
timestamp 1698431365
transform 1 0 1792 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_43
timestamp 1698431365
transform 1 0 6160 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_59
timestamp 1698431365
transform 1 0 7952 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_63
timestamp 1698431365
transform 1 0 8400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_74
timestamp 1698431365
transform 1 0 9632 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_78
timestamp 1698431365
transform 1 0 10080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_80
timestamp 1698431365
transform 1 0 10304 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_143
timestamp 1698431365
transform 1 0 17360 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_147
timestamp 1698431365
transform 1 0 17808 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_149
timestamp 1698431365
transform 1 0 18032 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_156
timestamp 1698431365
transform 1 0 18816 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_185
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_217
timestamp 1698431365
transform 1 0 25648 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_221
timestamp 1698431365
transform 1 0 26096 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_237
timestamp 1698431365
transform 1 0 27888 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_249
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_256
timestamp 1698431365
transform 1 0 30016 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_288
timestamp 1698431365
transform 1 0 33600 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_304
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_419
timestamp 1698431365
transform 1 0 48272 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_28
timestamp 1698431365
transform 1 0 4480 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_32
timestamp 1698431365
transform 1 0 4928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_36
timestamp 1698431365
transform 1 0 5376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_42
timestamp 1698431365
transform 1 0 6048 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_76
timestamp 1698431365
transform 1 0 9856 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_84
timestamp 1698431365
transform 1 0 10752 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_88
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_90
timestamp 1698431365
transform 1 0 11424 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_175
timestamp 1698431365
transform 1 0 20944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_179
timestamp 1698431365
transform 1 0 21392 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_195
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_221
timestamp 1698431365
transform 1 0 26096 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_229
timestamp 1698431365
transform 1 0 26992 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_246
timestamp 1698431365
transform 1 0 28896 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_250
timestamp 1698431365
transform 1 0 29344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_252
timestamp 1698431365
transform 1 0 29568 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_261
timestamp 1698431365
transform 1 0 30576 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_45
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_49
timestamp 1698431365
transform 1 0 6832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_62
timestamp 1698431365
transform 1 0 8288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_66
timestamp 1698431365
transform 1 0 8736 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_82
timestamp 1698431365
transform 1 0 10528 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_86
timestamp 1698431365
transform 1 0 10976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_88
timestamp 1698431365
transform 1 0 11200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_148
timestamp 1698431365
transform 1 0 17920 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_164
timestamp 1698431365
transform 1 0 19712 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_193
timestamp 1698431365
transform 1 0 22960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_195
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_215
timestamp 1698431365
transform 1 0 25424 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698431365
transform 1 0 27216 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698431365
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_267
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_271
timestamp 1698431365
transform 1 0 31696 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_287
timestamp 1698431365
transform 1 0 33488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_291
timestamp 1698431365
transform 1 0 33936 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_294
timestamp 1698431365
transform 1 0 34272 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_310
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_379
timestamp 1698431365
transform 1 0 43792 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_383
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_419
timestamp 1698431365
transform 1 0 48272 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_10
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_41
timestamp 1698431365
transform 1 0 5936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_45
timestamp 1698431365
transform 1 0 6384 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_61
timestamp 1698431365
transform 1 0 8176 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_127
timestamp 1698431365
transform 1 0 15568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_129
timestamp 1698431365
transform 1 0 15792 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_157
timestamp 1698431365
transform 1 0 18928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_163
timestamp 1698431365
transform 1 0 19600 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_172
timestamp 1698431365
transform 1 0 20608 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_180
timestamp 1698431365
transform 1 0 21504 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_184
timestamp 1698431365
transform 1 0 21952 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_186
timestamp 1698431365
transform 1 0 22176 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_189
timestamp 1698431365
transform 1 0 22512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_197
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_228
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_232
timestamp 1698431365
transform 1 0 27328 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_262
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698431365
transform 1 0 31136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_301
timestamp 1698431365
transform 1 0 35056 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_309
timestamp 1698431365
transform 1 0 35952 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_317
timestamp 1698431365
transform 1 0 36848 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_333
timestamp 1698431365
transform 1 0 38640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_337
timestamp 1698431365
transform 1 0 39088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_345
timestamp 1698431365
transform 1 0 39984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_51
timestamp 1698431365
transform 1 0 7056 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_83
timestamp 1698431365
transform 1 0 10640 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_99
timestamp 1698431365
transform 1 0 12432 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_132
timestamp 1698431365
transform 1 0 16128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_136
timestamp 1698431365
transform 1 0 16576 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_151
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_229
timestamp 1698431365
transform 1 0 26992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_233
timestamp 1698431365
transform 1 0 27440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_249
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_279
timestamp 1698431365
transform 1 0 32592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_305
timestamp 1698431365
transform 1 0 35504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_333
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_343
timestamp 1698431365
transform 1 0 39760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_347
timestamp 1698431365
transform 1 0 40208 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_379
timestamp 1698431365
transform 1 0 43792 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_383
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_403
timestamp 1698431365
transform 1 0 46480 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_411
timestamp 1698431365
transform 1 0 47376 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_28
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_52
timestamp 1698431365
transform 1 0 7168 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_56
timestamp 1698431365
transform 1 0 7616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_112
timestamp 1698431365
transform 1 0 13888 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_120
timestamp 1698431365
transform 1 0 14784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_122
timestamp 1698431365
transform 1 0 15008 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_131
timestamp 1698431365
transform 1 0 16016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_135
timestamp 1698431365
transform 1 0 16464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_154
timestamp 1698431365
transform 1 0 18592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_158
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_187
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_216
timestamp 1698431365
transform 1 0 25536 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_286
timestamp 1698431365
transform 1 0 33376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_306
timestamp 1698431365
transform 1 0 35616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_310
timestamp 1698431365
transform 1 0 36064 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_41
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_51
timestamp 1698431365
transform 1 0 7056 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_67
timestamp 1698431365
transform 1 0 8848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_89
timestamp 1698431365
transform 1 0 11312 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_93
timestamp 1698431365
transform 1 0 11760 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698431365
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698431365
transform 1 0 14000 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_164
timestamp 1698431365
transform 1 0 19712 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_168
timestamp 1698431365
transform 1 0 20160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698431365
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_207
timestamp 1698431365
transform 1 0 24528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_209
timestamp 1698431365
transform 1 0 24752 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_230
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_234
timestamp 1698431365
transform 1 0 27552 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_263
timestamp 1698431365
transform 1 0 30800 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_271
timestamp 1698431365
transform 1 0 31696 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_274
timestamp 1698431365
transform 1 0 32032 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_290
timestamp 1698431365
transform 1 0 33824 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_298
timestamp 1698431365
transform 1 0 34720 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_310
timestamp 1698431365
transform 1 0 36064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_364
timestamp 1698431365
transform 1 0 42112 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_380
timestamp 1698431365
transform 1 0 43904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_419
timestamp 1698431365
transform 1 0 48272 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_10
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_12
timestamp 1698431365
transform 1 0 2688 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_42
timestamp 1698431365
transform 1 0 6048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_46
timestamp 1698431365
transform 1 0 6496 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_54
timestamp 1698431365
transform 1 0 7392 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_91
timestamp 1698431365
transform 1 0 11536 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_107
timestamp 1698431365
transform 1 0 13328 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_111
timestamp 1698431365
transform 1 0 13776 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_167
timestamp 1698431365
transform 1 0 20048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_171
timestamp 1698431365
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_175
timestamp 1698431365
transform 1 0 20944 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_183
timestamp 1698431365
transform 1 0 21840 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_189
timestamp 1698431365
transform 1 0 22512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_199
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_203
timestamp 1698431365
transform 1 0 24080 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_207
timestamp 1698431365
transform 1 0 24528 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_241
timestamp 1698431365
transform 1 0 28336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_245
timestamp 1698431365
transform 1 0 28784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_253
timestamp 1698431365
transform 1 0 29680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_257
timestamp 1698431365
transform 1 0 30128 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_265
timestamp 1698431365
transform 1 0 31024 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_273
timestamp 1698431365
transform 1 0 31920 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_317
timestamp 1698431365
transform 1 0 36848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_321
timestamp 1698431365
transform 1 0 37296 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_329
timestamp 1698431365
transform 1 0 38192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_333
timestamp 1698431365
transform 1 0 38640 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_342
timestamp 1698431365
transform 1 0 39648 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_49
timestamp 1698431365
transform 1 0 6832 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_53
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_58
timestamp 1698431365
transform 1 0 7840 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_83
timestamp 1698431365
transform 1 0 10640 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_99
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_117
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_120
timestamp 1698431365
transform 1 0 14784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_124
timestamp 1698431365
transform 1 0 15232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_128
timestamp 1698431365
transform 1 0 15680 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_140
timestamp 1698431365
transform 1 0 17024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_144
timestamp 1698431365
transform 1 0 17472 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_148
timestamp 1698431365
transform 1 0 17920 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_209
timestamp 1698431365
transform 1 0 24752 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_217
timestamp 1698431365
transform 1 0 25648 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_221
timestamp 1698431365
transform 1 0 26096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_223
timestamp 1698431365
transform 1 0 26320 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_230
timestamp 1698431365
transform 1 0 27104 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_238
timestamp 1698431365
transform 1 0 28000 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_255
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_287
timestamp 1698431365
transform 1 0 33488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_295
timestamp 1698431365
transform 1 0 34384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_303
timestamp 1698431365
transform 1 0 35280 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_307
timestamp 1698431365
transform 1 0 35728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_333
timestamp 1698431365
transform 1 0 38640 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_343
timestamp 1698431365
transform 1 0 39760 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_375
timestamp 1698431365
transform 1 0 43344 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_419
timestamp 1698431365
transform 1 0 48272 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_104
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_108
timestamp 1698431365
transform 1 0 13440 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_127
timestamp 1698431365
transform 1 0 15568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_134
timestamp 1698431365
transform 1 0 16352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_138
timestamp 1698431365
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_144
timestamp 1698431365
transform 1 0 17472 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_147
timestamp 1698431365
transform 1 0 17808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_151
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_155
timestamp 1698431365
transform 1 0 18704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_168
timestamp 1698431365
transform 1 0 20160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_172
timestamp 1698431365
transform 1 0 20608 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_204
timestamp 1698431365
transform 1 0 24192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_228
timestamp 1698431365
transform 1 0 26880 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_232
timestamp 1698431365
transform 1 0 27328 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_262
timestamp 1698431365
transform 1 0 30688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_266
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_274
timestamp 1698431365
transform 1 0 32032 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_289
timestamp 1698431365
transform 1 0 33712 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_293
timestamp 1698431365
transform 1 0 34160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_295
timestamp 1698431365
transform 1 0 34384 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_303
timestamp 1698431365
transform 1 0 35280 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_335
timestamp 1698431365
transform 1 0 38864 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_343
timestamp 1698431365
transform 1 0 39760 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_347
timestamp 1698431365
transform 1 0 40208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_28
timestamp 1698431365
transform 1 0 4480 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_53
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_61
timestamp 1698431365
transform 1 0 8176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_77
timestamp 1698431365
transform 1 0 9968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_81
timestamp 1698431365
transform 1 0 10416 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_97
timestamp 1698431365
transform 1 0 12208 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_140
timestamp 1698431365
transform 1 0 17024 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_144
timestamp 1698431365
transform 1 0 17472 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_155
timestamp 1698431365
transform 1 0 18704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_157
timestamp 1698431365
transform 1 0 18928 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_179
timestamp 1698431365
transform 1 0 21392 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_218
timestamp 1698431365
transform 1 0 25760 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_222
timestamp 1698431365
transform 1 0 26208 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_238
timestamp 1698431365
transform 1 0 28000 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_293
timestamp 1698431365
transform 1 0 34160 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_297
timestamp 1698431365
transform 1 0 34608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_299
timestamp 1698431365
transform 1 0 34832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_310
timestamp 1698431365
transform 1 0 36064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_329
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_331
timestamp 1698431365
transform 1 0 38416 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_363
timestamp 1698431365
transform 1 0 42000 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_379
timestamp 1698431365
transform 1 0 43792 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_383
timestamp 1698431365
transform 1 0 44240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_51
timestamp 1698431365
transform 1 0 7056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_83
timestamp 1698431365
transform 1 0 10640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_87
timestamp 1698431365
transform 1 0 11088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_91
timestamp 1698431365
transform 1 0 11536 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_99
timestamp 1698431365
transform 1 0 12432 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_103
timestamp 1698431365
transform 1 0 12880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_105
timestamp 1698431365
transform 1 0 13104 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_129
timestamp 1698431365
transform 1 0 15792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_133
timestamp 1698431365
transform 1 0 16240 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698431365
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_146
timestamp 1698431365
transform 1 0 17696 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_189
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_193
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_197
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_205
timestamp 1698431365
transform 1 0 24304 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_208
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_248
timestamp 1698431365
transform 1 0 29120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_252
timestamp 1698431365
transform 1 0 29568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_268
timestamp 1698431365
transform 1 0 31360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_286
timestamp 1698431365
transform 1 0 33376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_288
timestamp 1698431365
transform 1 0 33600 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_321
timestamp 1698431365
transform 1 0 37296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_325
timestamp 1698431365
transform 1 0 37744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_329
timestamp 1698431365
transform 1 0 38192 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_358
timestamp 1698431365
transform 1 0 41440 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_362
timestamp 1698431365
transform 1 0 41888 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_379
timestamp 1698431365
transform 1 0 43792 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_411
timestamp 1698431365
transform 1 0 47376 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_33
timestamp 1698431365
transform 1 0 5040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_42
timestamp 1698431365
transform 1 0 6048 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_58
timestamp 1698431365
transform 1 0 7840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_60
timestamp 1698431365
transform 1 0 8064 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_82
timestamp 1698431365
transform 1 0 10528 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_86
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_88
timestamp 1698431365
transform 1 0 11200 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_111
timestamp 1698431365
transform 1 0 13776 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_119
timestamp 1698431365
transform 1 0 14672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_155
timestamp 1698431365
transform 1 0 18704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_168
timestamp 1698431365
transform 1 0 20160 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_172
timestamp 1698431365
transform 1 0 20608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_209
timestamp 1698431365
transform 1 0 24752 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_225
timestamp 1698431365
transform 1 0 26544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_229
timestamp 1698431365
transform 1 0 26992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_236
timestamp 1698431365
transform 1 0 27776 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_419
timestamp 1698431365
transform 1 0 48272 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_28
timestamp 1698431365
transform 1 0 4480 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_32
timestamp 1698431365
transform 1 0 4928 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_35
timestamp 1698431365
transform 1 0 5264 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_80
timestamp 1698431365
transform 1 0 10304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_92
timestamp 1698431365
transform 1 0 11648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_108
timestamp 1698431365
transform 1 0 13440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_118
timestamp 1698431365
transform 1 0 14560 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_134
timestamp 1698431365
transform 1 0 16352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_138
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_154
timestamp 1698431365
transform 1 0 18592 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_164
timestamp 1698431365
transform 1 0 19712 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_170
timestamp 1698431365
transform 1 0 20384 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_202
timestamp 1698431365
transform 1 0 23968 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_224
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_237
timestamp 1698431365
transform 1 0 27888 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_251
timestamp 1698431365
transform 1 0 29456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_255
timestamp 1698431365
transform 1 0 29904 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_271
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_290
timestamp 1698431365
transform 1 0 33824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_294
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_315
timestamp 1698431365
transform 1 0 36624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_319
timestamp 1698431365
transform 1 0 37072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698431365
transform 1 0 47936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_69
timestamp 1698431365
transform 1 0 9072 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_78
timestamp 1698431365
transform 1 0 10080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_82
timestamp 1698431365
transform 1 0 10528 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_98
timestamp 1698431365
transform 1 0 12320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_139
timestamp 1698431365
transform 1 0 16912 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_151
timestamp 1698431365
transform 1 0 18256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_155
timestamp 1698431365
transform 1 0 18704 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_189
timestamp 1698431365
transform 1 0 22512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_196
timestamp 1698431365
transform 1 0 23296 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_228
timestamp 1698431365
transform 1 0 26880 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_261
timestamp 1698431365
transform 1 0 30576 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_293
timestamp 1698431365
transform 1 0 34160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_295
timestamp 1698431365
transform 1 0 34384 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_356
timestamp 1698431365
transform 1 0 41216 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_372
timestamp 1698431365
transform 1 0 43008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_380
timestamp 1698431365
transform 1 0 43904 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_419
timestamp 1698431365
transform 1 0 48272 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_8
timestamp 1698431365
transform 1 0 2240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_12
timestamp 1698431365
transform 1 0 2688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_16
timestamp 1698431365
transform 1 0 3136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_26
timestamp 1698431365
transform 1 0 4256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_30
timestamp 1698431365
transform 1 0 4704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_34
timestamp 1698431365
transform 1 0 5152 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_90
timestamp 1698431365
transform 1 0 11424 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_102
timestamp 1698431365
transform 1 0 12768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_104
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_117
timestamp 1698431365
transform 1 0 14448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_133
timestamp 1698431365
transform 1 0 16240 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_150
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_152
timestamp 1698431365
transform 1 0 18368 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_164
timestamp 1698431365
transform 1 0 19712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_168
timestamp 1698431365
transform 1 0 20160 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_176
timestamp 1698431365
transform 1 0 21056 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_216
timestamp 1698431365
transform 1 0 25536 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_220
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_231
timestamp 1698431365
transform 1 0 27216 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_261
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_265
timestamp 1698431365
transform 1 0 31024 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_273
timestamp 1698431365
transform 1 0 31920 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_277
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_298
timestamp 1698431365
transform 1 0 34720 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_310
timestamp 1698431365
transform 1 0 36064 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_342
timestamp 1698431365
transform 1 0 39648 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_6
timestamp 1698431365
transform 1 0 2016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_43
timestamp 1698431365
transform 1 0 6160 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_56
timestamp 1698431365
transform 1 0 7616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_60
timestamp 1698431365
transform 1 0 8064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_64
timestamp 1698431365
transform 1 0 8512 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_77
timestamp 1698431365
transform 1 0 9968 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_93
timestamp 1698431365
transform 1 0 11760 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_95
timestamp 1698431365
transform 1 0 11984 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_157
timestamp 1698431365
transform 1 0 18928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_161
timestamp 1698431365
transform 1 0 19376 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_169
timestamp 1698431365
transform 1 0 20272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_187
timestamp 1698431365
transform 1 0 22288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_196
timestamp 1698431365
transform 1 0 23296 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_212
timestamp 1698431365
transform 1 0 25088 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_263
timestamp 1698431365
transform 1 0 30800 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_279
timestamp 1698431365
transform 1 0 32592 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_282
timestamp 1698431365
transform 1 0 32928 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_290
timestamp 1698431365
transform 1 0 33824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_294
timestamp 1698431365
transform 1 0 34272 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_296
timestamp 1698431365
transform 1 0 34496 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_303
timestamp 1698431365
transform 1 0 35280 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_307
timestamp 1698431365
transform 1 0 35728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_309
timestamp 1698431365
transform 1 0 35952 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_333
timestamp 1698431365
transform 1 0 38640 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_341
timestamp 1698431365
transform 1 0 39536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_362
timestamp 1698431365
transform 1 0 41888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_366
timestamp 1698431365
transform 1 0 42336 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_382
timestamp 1698431365
transform 1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_419
timestamp 1698431365
transform 1 0 48272 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_78
timestamp 1698431365
transform 1 0 10080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_83
timestamp 1698431365
transform 1 0 10640 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_91
timestamp 1698431365
transform 1 0 11536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_93
timestamp 1698431365
transform 1 0 11760 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_102
timestamp 1698431365
transform 1 0 12768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_110
timestamp 1698431365
transform 1 0 13664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_114
timestamp 1698431365
transform 1 0 14112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_118
timestamp 1698431365
transform 1 0 14560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_122
timestamp 1698431365
transform 1 0 15008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_126
timestamp 1698431365
transform 1 0 15456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_146
timestamp 1698431365
transform 1 0 17696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_148
timestamp 1698431365
transform 1 0 17920 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_162
timestamp 1698431365
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_166
timestamp 1698431365
transform 1 0 19936 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_174
timestamp 1698431365
transform 1 0 20832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_205
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_244
timestamp 1698431365
transform 1 0 28672 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_252
timestamp 1698431365
transform 1 0 29568 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_255
timestamp 1698431365
transform 1 0 29904 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_271
timestamp 1698431365
transform 1 0 31696 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_311
timestamp 1698431365
transform 1 0 36176 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_341
timestamp 1698431365
transform 1 0 39536 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_28
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_30
timestamp 1698431365
transform 1 0 4704 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_47
timestamp 1698431365
transform 1 0 6608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_51
timestamp 1698431365
transform 1 0 7056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_59
timestamp 1698431365
transform 1 0 7952 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_68
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_81
timestamp 1698431365
transform 1 0 10416 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_116
timestamp 1698431365
transform 1 0 14336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_118
timestamp 1698431365
transform 1 0 14560 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_129
timestamp 1698431365
transform 1 0 15792 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_163
timestamp 1698431365
transform 1 0 19600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_167
timestamp 1698431365
transform 1 0 20048 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_184
timestamp 1698431365
transform 1 0 21952 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_190
timestamp 1698431365
transform 1 0 22624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_194
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_226
timestamp 1698431365
transform 1 0 26656 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_242
timestamp 1698431365
transform 1 0 28448 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_297
timestamp 1698431365
transform 1 0 34608 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_349
timestamp 1698431365
transform 1 0 40432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_351
timestamp 1698431365
transform 1 0 40656 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_358
timestamp 1698431365
transform 1 0 41440 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_374
timestamp 1698431365
transform 1 0 43232 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_382
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_384
timestamp 1698431365
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_403
timestamp 1698431365
transform 1 0 46480 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_411
timestamp 1698431365
transform 1 0 47376 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_6
timestamp 1698431365
transform 1 0 2016 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_36
timestamp 1698431365
transform 1 0 5376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_40
timestamp 1698431365
transform 1 0 5824 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_48
timestamp 1698431365
transform 1 0 6720 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_52
timestamp 1698431365
transform 1 0 7168 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_54
timestamp 1698431365
transform 1 0 7392 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_61
timestamp 1698431365
transform 1 0 8176 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_97
timestamp 1698431365
transform 1 0 12208 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_104
timestamp 1698431365
transform 1 0 12992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_108
timestamp 1698431365
transform 1 0 13440 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_134
timestamp 1698431365
transform 1 0 16352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_165
timestamp 1698431365
transform 1 0 19824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_169
timestamp 1698431365
transform 1 0 20272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_173
timestamp 1698431365
transform 1 0 20720 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698431365
transform 1 0 24304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_228
timestamp 1698431365
transform 1 0 26880 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_230
timestamp 1698431365
transform 1 0 27104 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_248
timestamp 1698431365
transform 1 0 29120 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_252
timestamp 1698431365
transform 1 0 29568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_256
timestamp 1698431365
transform 1 0 30016 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_272
timestamp 1698431365
transform 1 0 31808 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_297
timestamp 1698431365
transform 1 0 34608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_301
timestamp 1698431365
transform 1 0 35056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_305
timestamp 1698431365
transform 1 0 35504 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_337
timestamp 1698431365
transform 1 0 39088 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_345
timestamp 1698431365
transform 1 0 39984 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_10
timestamp 1698431365
transform 1 0 2464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_55
timestamp 1698431365
transform 1 0 7504 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_62
timestamp 1698431365
transform 1 0 8288 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_70
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_74
timestamp 1698431365
transform 1 0 9632 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_85
timestamp 1698431365
transform 1 0 10864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_89
timestamp 1698431365
transform 1 0 11312 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_97
timestamp 1698431365
transform 1 0 12208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_115
timestamp 1698431365
transform 1 0 14224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_167
timestamp 1698431365
transform 1 0 20048 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_192
timestamp 1698431365
transform 1 0 22848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_199
timestamp 1698431365
transform 1 0 23632 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_231
timestamp 1698431365
transform 1 0 27216 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_239
timestamp 1698431365
transform 1 0 28112 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_243
timestamp 1698431365
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_253
timestamp 1698431365
transform 1 0 29680 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_285
timestamp 1698431365
transform 1 0 33264 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_301
timestamp 1698431365
transform 1 0 35056 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_309
timestamp 1698431365
transform 1 0 35952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_349
timestamp 1698431365
transform 1 0 40432 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_353
timestamp 1698431365
transform 1 0 40880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_357
timestamp 1698431365
transform 1 0 41328 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_373
timestamp 1698431365
transform 1 0 43120 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_419
timestamp 1698431365
transform 1 0 48272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_28
timestamp 1698431365
transform 1 0 4480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_32
timestamp 1698431365
transform 1 0 4928 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_62
timestamp 1698431365
transform 1 0 8288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_84
timestamp 1698431365
transform 1 0 10752 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_88
timestamp 1698431365
transform 1 0 11200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_104
timestamp 1698431365
transform 1 0 12992 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_110
timestamp 1698431365
transform 1 0 13664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_114
timestamp 1698431365
transform 1 0 14112 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_150
timestamp 1698431365
transform 1 0 18144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_157
timestamp 1698431365
transform 1 0 18928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_161
timestamp 1698431365
transform 1 0 19376 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_177
timestamp 1698431365
transform 1 0 21168 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_216
timestamp 1698431365
transform 1 0 25536 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_224
timestamp 1698431365
transform 1 0 26432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_246
timestamp 1698431365
transform 1 0 28896 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_254
timestamp 1698431365
transform 1 0 29792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_256
timestamp 1698431365
transform 1 0 30016 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_272
timestamp 1698431365
transform 1 0 31808 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_286
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_288
timestamp 1698431365
transform 1 0 33600 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_304
timestamp 1698431365
transform 1 0 35392 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_308
timestamp 1698431365
transform 1 0 35840 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_312
timestamp 1698431365
transform 1 0 36288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_316
timestamp 1698431365
transform 1 0 36736 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_348
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698431365
transform 1 0 47936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_45
timestamp 1698431365
transform 1 0 6384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_55
timestamp 1698431365
transform 1 0 7504 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_87
timestamp 1698431365
transform 1 0 11088 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_103
timestamp 1698431365
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_126
timestamp 1698431365
transform 1 0 15456 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_130
timestamp 1698431365
transform 1 0 15904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_134
timestamp 1698431365
transform 1 0 16352 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_140
timestamp 1698431365
transform 1 0 17024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_144
timestamp 1698431365
transform 1 0 17472 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_148
timestamp 1698431365
transform 1 0 17920 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_164
timestamp 1698431365
transform 1 0 19712 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_172
timestamp 1698431365
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_189
timestamp 1698431365
transform 1 0 22512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_193
timestamp 1698431365
transform 1 0 22960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_195
timestamp 1698431365
transform 1 0 23184 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_204
timestamp 1698431365
transform 1 0 24192 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_220
timestamp 1698431365
transform 1 0 25984 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_228
timestamp 1698431365
transform 1 0 26880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_235
timestamp 1698431365
transform 1 0 27664 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_307
timestamp 1698431365
transform 1 0 35728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_337
timestamp 1698431365
transform 1 0 39088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_345
timestamp 1698431365
transform 1 0 39984 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_377
timestamp 1698431365
transform 1 0 43568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_419
timestamp 1698431365
transform 1 0 48272 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_28
timestamp 1698431365
transform 1 0 4480 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_44
timestamp 1698431365
transform 1 0 6272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_46
timestamp 1698431365
transform 1 0 6496 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_53
timestamp 1698431365
transform 1 0 7280 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_88
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_96
timestamp 1698431365
transform 1 0 12096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_100
timestamp 1698431365
transform 1 0 12544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_102
timestamp 1698431365
transform 1 0 12768 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_114
timestamp 1698431365
transform 1 0 14112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_118
timestamp 1698431365
transform 1 0 14560 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_134
timestamp 1698431365
transform 1 0 16352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_138
timestamp 1698431365
transform 1 0 16800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_158
timestamp 1698431365
transform 1 0 19040 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_166
timestamp 1698431365
transform 1 0 19936 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_168
timestamp 1698431365
transform 1 0 20160 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_175
timestamp 1698431365
transform 1 0 20944 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1698431365
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_224
timestamp 1698431365
transform 1 0 26432 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_242
timestamp 1698431365
transform 1 0 28448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_246
timestamp 1698431365
transform 1 0 28896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_250
timestamp 1698431365
transform 1 0 29344 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_266
timestamp 1698431365
transform 1 0 31136 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_274
timestamp 1698431365
transform 1 0 32032 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_33
timestamp 1698431365
transform 1 0 5040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_41
timestamp 1698431365
transform 1 0 5936 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_51
timestamp 1698431365
transform 1 0 7056 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_65
timestamp 1698431365
transform 1 0 8624 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_69
timestamp 1698431365
transform 1 0 9072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_72
timestamp 1698431365
transform 1 0 9408 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_88
timestamp 1698431365
transform 1 0 11200 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_102
timestamp 1698431365
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_111
timestamp 1698431365
transform 1 0 13776 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_143
timestamp 1698431365
transform 1 0 17360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_157
timestamp 1698431365
transform 1 0 18928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_161
timestamp 1698431365
transform 1 0 19376 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_165
timestamp 1698431365
transform 1 0 19824 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_185
timestamp 1698431365
transform 1 0 22064 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_198
timestamp 1698431365
transform 1 0 23520 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_202
timestamp 1698431365
transform 1 0 23968 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_218
timestamp 1698431365
transform 1 0 25760 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_226
timestamp 1698431365
transform 1 0 26656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_230
timestamp 1698431365
transform 1 0 27104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_232
timestamp 1698431365
transform 1 0 27328 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_403
timestamp 1698431365
transform 1 0 46480 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_411
timestamp 1698431365
transform 1 0 47376 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_74
timestamp 1698431365
transform 1 0 9632 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_96
timestamp 1698431365
transform 1 0 12096 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_128
timestamp 1698431365
transform 1 0 15680 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_155
timestamp 1698431365
transform 1 0 18704 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_171
timestamp 1698431365
transform 1 0 20496 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_179
timestamp 1698431365
transform 1 0 21392 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_183
timestamp 1698431365
transform 1 0 21840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_190
timestamp 1698431365
transform 1 0 22624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_194
timestamp 1698431365
transform 1 0 23072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_203
timestamp 1698431365
transform 1 0 24080 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_207
timestamp 1698431365
transform 1 0 24528 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_228
timestamp 1698431365
transform 1 0 26880 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_232
timestamp 1698431365
transform 1 0 27328 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_234
timestamp 1698431365
transform 1 0 27552 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_264
timestamp 1698431365
transform 1 0 30912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_268
timestamp 1698431365
transform 1 0 31360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_53
timestamp 1698431365
transform 1 0 7280 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_55
timestamp 1698431365
transform 1 0 7504 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_62
timestamp 1698431365
transform 1 0 8288 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_68
timestamp 1698431365
transform 1 0 8960 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_72
timestamp 1698431365
transform 1 0 9408 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_103
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_111
timestamp 1698431365
transform 1 0 13776 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_119
timestamp 1698431365
transform 1 0 14672 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_158
timestamp 1698431365
transform 1 0 19040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_162
timestamp 1698431365
transform 1 0 19488 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_168
timestamp 1698431365
transform 1 0 20160 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_186
timestamp 1698431365
transform 1 0 22176 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_195
timestamp 1698431365
transform 1 0 23184 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_207
timestamp 1698431365
transform 1 0 24528 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_211
timestamp 1698431365
transform 1 0 24976 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_227
timestamp 1698431365
transform 1 0 26768 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_235
timestamp 1698431365
transform 1 0 27664 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_239
timestamp 1698431365
transform 1 0 28112 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_251
timestamp 1698431365
transform 1 0 29456 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_333
timestamp 1698431365
transform 1 0 38640 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_341
timestamp 1698431365
transform 1 0 39536 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_344
timestamp 1698431365
transform 1 0 39872 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_348
timestamp 1698431365
transform 1 0 40320 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_365
timestamp 1698431365
transform 1 0 42224 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_391
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_393
timestamp 1698431365
transform 1 0 45360 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_28
timestamp 1698431365
transform 1 0 4480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_32
timestamp 1698431365
transform 1 0 4928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_36
timestamp 1698431365
transform 1 0 5376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_40
timestamp 1698431365
transform 1 0 5824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_44
timestamp 1698431365
transform 1 0 6272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_46
timestamp 1698431365
transform 1 0 6496 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_57
timestamp 1698431365
transform 1 0 7728 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_63
timestamp 1698431365
transform 1 0 8400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_67
timestamp 1698431365
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_85
timestamp 1698431365
transform 1 0 10864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_87
timestamp 1698431365
transform 1 0 11088 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_117
timestamp 1698431365
transform 1 0 14448 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_121
timestamp 1698431365
transform 1 0 14896 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_137
timestamp 1698431365
transform 1 0 16688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698431365
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_151
timestamp 1698431365
transform 1 0 18256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_155
timestamp 1698431365
transform 1 0 18704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_157
timestamp 1698431365
transform 1 0 18928 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_166
timestamp 1698431365
transform 1 0 19936 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_168
timestamp 1698431365
transform 1 0 20160 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_241
timestamp 1698431365
transform 1 0 28336 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_245
timestamp 1698431365
transform 1 0 28784 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_260
timestamp 1698431365
transform 1 0 30464 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_264
timestamp 1698431365
transform 1 0 30912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_272
timestamp 1698431365
transform 1 0 31808 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_288
timestamp 1698431365
transform 1 0 33600 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_320
timestamp 1698431365
transform 1 0 37184 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_336
timestamp 1698431365
transform 1 0 38976 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_344
timestamp 1698431365
transform 1 0 39872 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698431365
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_384
timestamp 1698431365
transform 1 0 44352 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_33
timestamp 1698431365
transform 1 0 5040 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_39
timestamp 1698431365
transform 1 0 5712 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_69
timestamp 1698431365
transform 1 0 9072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_73
timestamp 1698431365
transform 1 0 9520 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_81
timestamp 1698431365
transform 1 0 10416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_85
timestamp 1698431365
transform 1 0 10864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_87
timestamp 1698431365
transform 1 0 11088 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_94
timestamp 1698431365
transform 1 0 11872 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_102
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_115
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_117
timestamp 1698431365
transform 1 0 14448 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_126
timestamp 1698431365
transform 1 0 15456 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_130
timestamp 1698431365
transform 1 0 15904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_132
timestamp 1698431365
transform 1 0 16128 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_162
timestamp 1698431365
transform 1 0 19488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_166
timestamp 1698431365
transform 1 0 19936 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_181
timestamp 1698431365
transform 1 0 21616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_193
timestamp 1698431365
transform 1 0 22960 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_197
timestamp 1698431365
transform 1 0 23408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_231
timestamp 1698431365
transform 1 0 27216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_297
timestamp 1698431365
transform 1 0 34608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_301
timestamp 1698431365
transform 1 0 35056 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_308
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698431365
transform 1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_413
timestamp 1698431365
transform 1 0 47600 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_417
timestamp 1698431365
transform 1 0 48048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_419
timestamp 1698431365
transform 1 0 48272 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_60
timestamp 1698431365
transform 1 0 8064 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_67
timestamp 1698431365
transform 1 0 8848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_69
timestamp 1698431365
transform 1 0 9072 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_84
timestamp 1698431365
transform 1 0 10752 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_88
timestamp 1698431365
transform 1 0 11200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_90
timestamp 1698431365
transform 1 0 11424 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_97
timestamp 1698431365
transform 1 0 12208 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_101
timestamp 1698431365
transform 1 0 12656 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_104
timestamp 1698431365
transform 1 0 12992 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_146
timestamp 1698431365
transform 1 0 17696 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_178
timestamp 1698431365
transform 1 0 21280 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_181
timestamp 1698431365
transform 1 0 21616 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_197
timestamp 1698431365
transform 1 0 23408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_205
timestamp 1698431365
transform 1 0 24304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_214
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_221
timestamp 1698431365
transform 1 0 26096 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_255
timestamp 1698431365
transform 1 0 29904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_259
timestamp 1698431365
transform 1 0 30352 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_267
timestamp 1698431365
transform 1 0 31248 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_274
timestamp 1698431365
transform 1 0 32032 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_278
timestamp 1698431365
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_334
timestamp 1698431365
transform 1 0 38752 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_404
timestamp 1698431365
transform 1 0 46592 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_36
timestamp 1698431365
transform 1 0 5376 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_45
timestamp 1698431365
transform 1 0 6384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_49
timestamp 1698431365
transform 1 0 6832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_51
timestamp 1698431365
transform 1 0 7056 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_54
timestamp 1698431365
transform 1 0 7392 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_58
timestamp 1698431365
transform 1 0 7840 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_61
timestamp 1698431365
transform 1 0 8176 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_70
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_72
timestamp 1698431365
transform 1 0 9408 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_79
timestamp 1698431365
transform 1 0 10192 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_91
timestamp 1698431365
transform 1 0 11536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_95
timestamp 1698431365
transform 1 0 11984 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_106
timestamp 1698431365
transform 1 0 13216 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_115
timestamp 1698431365
transform 1 0 14224 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_127
timestamp 1698431365
transform 1 0 15568 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_131
timestamp 1698431365
transform 1 0 16016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_133
timestamp 1698431365
transform 1 0 16240 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_144
timestamp 1698431365
transform 1 0 17472 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_151
timestamp 1698431365
transform 1 0 18256 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_163
timestamp 1698431365
transform 1 0 19600 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_167
timestamp 1698431365
transform 1 0 20048 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_178
timestamp 1698431365
transform 1 0 21280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_180
timestamp 1698431365
transform 1 0 21504 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_187
timestamp 1698431365
transform 1 0 22288 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_199
timestamp 1698431365
transform 1 0 23632 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_203
timestamp 1698431365
transform 1 0 24080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_206
timestamp 1698431365
transform 1 0 24416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_210
timestamp 1698431365
transform 1 0 24864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_240
timestamp 1698431365
transform 1 0 28224 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_267
timestamp 1698431365
transform 1 0 31248 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_271
timestamp 1698431365
transform 1 0 31696 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_300
timestamp 1698431365
transform 1 0 34944 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_304
timestamp 1698431365
transform 1 0 35392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_334
timestamp 1698431365
transform 1 0 38752 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_338
timestamp 1698431365
transform 1 0 39200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_368
timestamp 1698431365
transform 1 0 42560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_372
timestamp 1698431365
transform 1 0 43008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_402
timestamp 1698431365
transform 1 0 46368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_406
timestamp 1698431365
transform 1 0 46816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_410
timestamp 1698431365
transform 1 0 47264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  hold1
timestamp 1698431365
transform -1 0 12208 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold2
timestamp 1698431365
transform -1 0 8176 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold3
timestamp 1698431365
transform -1 0 7280 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold4
timestamp 1698431365
transform -1 0 8288 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold5
timestamp 1698431365
transform -1 0 7280 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold6
timestamp 1698431365
transform -1 0 8960 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  hold7
timestamp 1698431365
transform -1 0 11872 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold8
timestamp 1698431365
transform -1 0 8288 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 48384 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 48384 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 48384 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 48384 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 36512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input11
timestamp 1698431365
transform -1 0 37744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input13
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input14
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input15
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input16
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input17
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input20
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input21
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 17584 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 19600 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 21280 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 22288 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 23632 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 4480 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 4480 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 7392 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 8176 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 9520 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 10864 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input33
timestamp 1698431365
transform 1 0 12096 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input34
timestamp 1698431365
transform 1 0 13552 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 14896 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform -1 0 48384 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform -1 0 48384 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform -1 0 48384 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input39
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input40
timestamp 1698431365
transform -1 0 48384 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input41
timestamp 1698431365
transform -1 0 48384 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output42 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4480 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output43
timestamp 1698431365
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output44
timestamp 1698431365
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output45
timestamp 1698431365
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output46
timestamp 1698431365
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output47
timestamp 1698431365
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output48
timestamp 1698431365
transform -1 0 4480 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49
timestamp 1698431365
transform -1 0 4480 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698431365
transform -1 0 4480 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698431365
transform -1 0 27888 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698431365
transform 1 0 26992 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698431365
transform 1 0 28896 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698431365
transform 1 0 33040 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output58
timestamp 1698431365
transform -1 0 7728 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output59
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output60
timestamp 1698431365
transform -1 0 12320 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output61
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output62
timestamp 1698431365
transform 1 0 12880 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output63
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output64
timestamp 1698431365
transform -1 0 19824 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output65
timestamp 1698431365
transform -1 0 21840 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output66
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output67
timestamp 1698431365
transform 1 0 24304 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output68
timestamp 1698431365
transform 1 0 39648 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output69
timestamp 1698431365
transform 1 0 39760 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output70
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output71
timestamp 1698431365
transform 1 0 43456 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output72
timestamp 1698431365
transform 1 0 43680 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output73
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output74
timestamp 1698431365
transform 1 0 25088 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output75
timestamp 1698431365
transform 1 0 26992 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output76
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output77
timestamp 1698431365
transform 1 0 29680 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output78
timestamp 1698431365
transform 1 0 32032 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output79
timestamp 1698431365
transform -1 0 35840 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output80
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output81
timestamp 1698431365
transform 1 0 35840 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output82
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83
timestamp 1698431365
transform -1 0 42560 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84
timestamp 1698431365
transform 1 0 41104 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform -1 0 46368 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform -1 0 4480 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform -1 0 4480 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform -1 0 4480 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform -1 0 4480 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform -1 0 4480 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform -1 0 4480 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92
timestamp 1698431365
transform -1 0 4480 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform -1 0 7392 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform 1 0 45472 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform 1 0 45472 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_123
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_125
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_126
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_128
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_129
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_130
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_132
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_134
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_135
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_136
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_137
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_144
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_145
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_150
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_151
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_152
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_155
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_156
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_157
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_158
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_159
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_161
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_162
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_163
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_164
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_165
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_166
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_167
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_168
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_169
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_170
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_172
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_173
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_174
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_175
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_177
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_178
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_185
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_186
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_187
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_188
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_189
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_190
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_191
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_192
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_194
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_195
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_196
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_197
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_198
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_199
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_200
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_201
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_202
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_203
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_205
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_206
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_207
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_208
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_209
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_210
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_211
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_212
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_213
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_214
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_216
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_217
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_218
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_219
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_220
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_221
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_222
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_223
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_224
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_225
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_227
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_228
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_229
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_230
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_231
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_232
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_233
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_234
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_235
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_236
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_238
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_239
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_240
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_241
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_242
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_243
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_244
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_245
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_246
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_247
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_249
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_250
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_251
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_252
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_253
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_254
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_255
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_256
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_257
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_258
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_260
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_261
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_262
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_263
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_264
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_265
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_266
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_267
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_268
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_269
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_271
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_272
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_273
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_274
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_275
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_276
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_277
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_278
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_279
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_280
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_282
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_283
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_284
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_285
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_286
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_287
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_288
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_289
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_290
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_291
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_293
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_294
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_295
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_296
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_297
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_298
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_299
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_300
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_301
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_302
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_304
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_305
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_306
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_307
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_308
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_309
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_310
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_311
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_312
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_313
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_315
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_316
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_317
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_318
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_319
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_320
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_321
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_322
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_323
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_324
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_326
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_327
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_328
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_329
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_330
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_331
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_332
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_333
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_334
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_335
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_337
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_338
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_339
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_340
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_341
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_342
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_343
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_344
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_345
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_346
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_348
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_349
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_350
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_351
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_352
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_353
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_354
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_355
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_356
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_357
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_359
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_360
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_361
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_362
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_363
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_364
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_365
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_366
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_367
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_368
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_370
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_371
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_372
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_373
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_374
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_375
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_376
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_377
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_378
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_379
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_381
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_382
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_383
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_384
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_385
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_386
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_387
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_388
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_389
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_390
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_392
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_393
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_394
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_395
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_396
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_397
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_398
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_399
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_400
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_401
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_408
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_409
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_410
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_411
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_412
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_413
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_414
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_415
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_416
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_417
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_418
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_419
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_420
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_421
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_422
timestamp 1698431365
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_423
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_424
timestamp 1698431365
transform 1 0 47040 0 1 45472
box -86 -86 310 870
<< labels >>
flabel metal3 s 49200 30240 50000 30352 0 FreeSans 448 0 0 0 DAC_clk
port 0 nsew signal input
flabel metal3 s 49200 35616 50000 35728 0 FreeSans 448 0 0 0 DAC_d1
port 1 nsew signal input
flabel metal3 s 49200 40992 50000 41104 0 FreeSans 448 0 0 0 DAC_d2
port 2 nsew signal input
flabel metal3 s 49200 46368 50000 46480 0 FreeSans 448 0 0 0 DAC_le
port 3 nsew signal input
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 RXD
port 4 nsew signal tristate
flabel metal3 s 0 33376 800 33488 0 FreeSans 448 0 0 0 TXD
port 5 nsew signal input
flabel metal3 s 0 2016 800 2128 0 FreeSans 448 0 0 0 addr[0]
port 6 nsew signal input
flabel metal3 s 0 3584 800 3696 0 FreeSans 448 0 0 0 addr[1]
port 7 nsew signal input
flabel metal3 s 0 5152 800 5264 0 FreeSans 448 0 0 0 addr[2]
port 8 nsew signal input
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 addr[3]
port 9 nsew signal input
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 bus_cyc
port 10 nsew signal input
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 bus_we
port 11 nsew signal input
flabel metal3 s 0 8288 800 8400 0 FreeSans 448 0 0 0 data_in[0]
port 12 nsew signal input
flabel metal3 s 0 9856 800 9968 0 FreeSans 448 0 0 0 data_in[1]
port 13 nsew signal input
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 data_in[2]
port 14 nsew signal input
flabel metal3 s 0 12992 800 13104 0 FreeSans 448 0 0 0 data_in[3]
port 15 nsew signal input
flabel metal3 s 0 14560 800 14672 0 FreeSans 448 0 0 0 data_in[4]
port 16 nsew signal input
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 data_in[5]
port 17 nsew signal input
flabel metal3 s 0 17696 800 17808 0 FreeSans 448 0 0 0 data_in[6]
port 18 nsew signal input
flabel metal3 s 0 19264 800 19376 0 FreeSans 448 0 0 0 data_in[7]
port 19 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 data_out[0]
port 20 nsew signal tristate
flabel metal3 s 0 22400 800 22512 0 FreeSans 448 0 0 0 data_out[1]
port 21 nsew signal tristate
flabel metal3 s 0 23968 800 24080 0 FreeSans 448 0 0 0 data_out[2]
port 22 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 data_out[3]
port 23 nsew signal tristate
flabel metal3 s 0 27104 800 27216 0 FreeSans 448 0 0 0 data_out[4]
port 24 nsew signal tristate
flabel metal3 s 0 28672 800 28784 0 FreeSans 448 0 0 0 data_out[5]
port 25 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 data_out[6]
port 26 nsew signal tristate
flabel metal3 s 0 31808 800 31920 0 FreeSans 448 0 0 0 data_out[7]
port 27 nsew signal tristate
flabel metal2 s 2688 49200 2800 50000 0 FreeSans 448 90 0 0 io_in[0]
port 28 nsew signal input
flabel metal2 s 16128 49200 16240 50000 0 FreeSans 448 90 0 0 io_in[10]
port 29 nsew signal input
flabel metal2 s 17472 49200 17584 50000 0 FreeSans 448 90 0 0 io_in[11]
port 30 nsew signal input
flabel metal2 s 18816 49200 18928 50000 0 FreeSans 448 90 0 0 io_in[12]
port 31 nsew signal input
flabel metal2 s 20160 49200 20272 50000 0 FreeSans 448 90 0 0 io_in[13]
port 32 nsew signal input
flabel metal2 s 21504 49200 21616 50000 0 FreeSans 448 90 0 0 io_in[14]
port 33 nsew signal input
flabel metal2 s 22848 49200 22960 50000 0 FreeSans 448 90 0 0 io_in[15]
port 34 nsew signal input
flabel metal2 s 4032 49200 4144 50000 0 FreeSans 448 90 0 0 io_in[1]
port 35 nsew signal input
flabel metal2 s 5376 49200 5488 50000 0 FreeSans 448 90 0 0 io_in[2]
port 36 nsew signal input
flabel metal2 s 6720 49200 6832 50000 0 FreeSans 448 90 0 0 io_in[3]
port 37 nsew signal input
flabel metal2 s 8064 49200 8176 50000 0 FreeSans 448 90 0 0 io_in[4]
port 38 nsew signal input
flabel metal2 s 9408 49200 9520 50000 0 FreeSans 448 90 0 0 io_in[5]
port 39 nsew signal input
flabel metal2 s 10752 49200 10864 50000 0 FreeSans 448 90 0 0 io_in[6]
port 40 nsew signal input
flabel metal2 s 12096 49200 12208 50000 0 FreeSans 448 90 0 0 io_in[7]
port 41 nsew signal input
flabel metal2 s 13440 49200 13552 50000 0 FreeSans 448 90 0 0 io_in[8]
port 42 nsew signal input
flabel metal2 s 14784 49200 14896 50000 0 FreeSans 448 90 0 0 io_in[9]
port 43 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 44 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 io_oeb[10]
port 45 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 io_oeb[11]
port 46 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 io_oeb[12]
port 47 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 io_oeb[13]
port 48 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 io_oeb[14]
port 49 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 io_oeb[15]
port 50 nsew signal tristate
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 51 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 io_oeb[2]
port 52 nsew signal tristate
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 53 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 io_oeb[4]
port 54 nsew signal tristate
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 io_oeb[5]
port 55 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 io_oeb[6]
port 56 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 io_oeb[7]
port 57 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 58 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 59 nsew signal tristate
flabel metal2 s 24192 49200 24304 50000 0 FreeSans 448 90 0 0 io_out[0]
port 60 nsew signal tristate
flabel metal2 s 37632 49200 37744 50000 0 FreeSans 448 90 0 0 io_out[10]
port 61 nsew signal tristate
flabel metal2 s 38976 49200 39088 50000 0 FreeSans 448 90 0 0 io_out[11]
port 62 nsew signal tristate
flabel metal2 s 40320 49200 40432 50000 0 FreeSans 448 90 0 0 io_out[12]
port 63 nsew signal tristate
flabel metal2 s 41664 49200 41776 50000 0 FreeSans 448 90 0 0 io_out[13]
port 64 nsew signal tristate
flabel metal2 s 43008 49200 43120 50000 0 FreeSans 448 90 0 0 io_out[14]
port 65 nsew signal tristate
flabel metal2 s 44352 49200 44464 50000 0 FreeSans 448 90 0 0 io_out[15]
port 66 nsew signal tristate
flabel metal2 s 25536 49200 25648 50000 0 FreeSans 448 90 0 0 io_out[1]
port 67 nsew signal tristate
flabel metal2 s 26880 49200 26992 50000 0 FreeSans 448 90 0 0 io_out[2]
port 68 nsew signal tristate
flabel metal2 s 28224 49200 28336 50000 0 FreeSans 448 90 0 0 io_out[3]
port 69 nsew signal tristate
flabel metal2 s 29568 49200 29680 50000 0 FreeSans 448 90 0 0 io_out[4]
port 70 nsew signal tristate
flabel metal2 s 30912 49200 31024 50000 0 FreeSans 448 90 0 0 io_out[5]
port 71 nsew signal tristate
flabel metal2 s 32256 49200 32368 50000 0 FreeSans 448 90 0 0 io_out[6]
port 72 nsew signal tristate
flabel metal2 s 33600 49200 33712 50000 0 FreeSans 448 90 0 0 io_out[7]
port 73 nsew signal tristate
flabel metal2 s 34944 49200 35056 50000 0 FreeSans 448 90 0 0 io_out[8]
port 74 nsew signal tristate
flabel metal2 s 36288 49200 36400 50000 0 FreeSans 448 90 0 0 io_out[9]
port 75 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 irq0
port 76 nsew signal tristate
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 irq6
port 77 nsew signal tristate
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 irq7
port 78 nsew signal tristate
flabel metal3 s 0 36512 800 36624 0 FreeSans 448 0 0 0 la_data_out[0]
port 79 nsew signal tristate
flabel metal3 s 0 38080 800 38192 0 FreeSans 448 0 0 0 la_data_out[1]
port 80 nsew signal tristate
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 la_data_out[2]
port 81 nsew signal tristate
flabel metal3 s 0 41216 800 41328 0 FreeSans 448 0 0 0 la_data_out[3]
port 82 nsew signal tristate
flabel metal3 s 0 42784 800 42896 0 FreeSans 448 0 0 0 la_data_out[4]
port 83 nsew signal tristate
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 la_data_out[5]
port 84 nsew signal tristate
flabel metal3 s 0 45920 800 46032 0 FreeSans 448 0 0 0 la_data_out[6]
port 85 nsew signal tristate
flabel metal3 s 0 47488 800 47600 0 FreeSans 448 0 0 0 la_data_out[7]
port 86 nsew signal tristate
flabel metal3 s 49200 14112 50000 14224 0 FreeSans 448 0 0 0 pwm0
port 87 nsew signal input
flabel metal3 s 49200 19488 50000 19600 0 FreeSans 448 0 0 0 pwm1
port 88 nsew signal input
flabel metal3 s 49200 24864 50000 24976 0 FreeSans 448 0 0 0 pwm2
port 89 nsew signal input
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 rst
port 90 nsew signal input
flabel metal2 s 45696 49200 45808 50000 0 FreeSans 448 90 0 0 tmr0_clk
port 91 nsew signal tristate
flabel metal3 s 49200 3360 50000 3472 0 FreeSans 448 0 0 0 tmr0_o
port 92 nsew signal input
flabel metal2 s 47040 49200 47152 50000 0 FreeSans 448 90 0 0 tmr1_clk
port 93 nsew signal tristate
flabel metal3 s 49200 8736 50000 8848 0 FreeSans 448 0 0 0 tmr1_o
port 94 nsew signal input
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 95 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 95 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 96 nsew ground bidirectional
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 wb_clk_i
port 97 nsew signal input
rlabel metal1 24976 46256 24976 46256 0 vdd
rlabel metal1 24976 45472 24976 45472 0 vss
rlabel metal2 48216 30632 48216 30632 0 DAC_clk
rlabel metal2 48216 36008 48216 36008 0 DAC_d1
rlabel metal3 48762 41048 48762 41048 0 DAC_d2
rlabel metal2 48216 46144 48216 46144 0 DAC_le
rlabel metal2 13272 30632 13272 30632 0 DDRA\[0\]
rlabel metal2 6664 20272 6664 20272 0 DDRA\[1\]
rlabel metal2 8008 18312 8008 18312 0 DDRA\[2\]
rlabel metal2 6104 11872 6104 11872 0 DDRA\[3\]
rlabel metal2 11648 9912 11648 9912 0 DDRA\[4\]
rlabel metal2 15512 9352 15512 9352 0 DDRA\[5\]
rlabel metal2 14840 11536 14840 11536 0 DDRA\[6\]
rlabel metal3 16968 25816 16968 25816 0 DDRA\[7\]
rlabel metal2 20328 21280 20328 21280 0 DDRB\[0\]
rlabel metal2 9912 11592 9912 11592 0 DDRB\[1\]
rlabel metal2 23016 6160 23016 6160 0 DDRB\[2\]
rlabel metal2 24696 23408 24696 23408 0 DDRB\[3\]
rlabel metal2 25928 9352 25928 9352 0 DDRB\[4\]
rlabel metal2 27272 14056 27272 14056 0 DDRB\[5\]
rlabel metal3 19152 17080 19152 17080 0 DDRB\[6\]
rlabel metal2 19376 19096 19376 19096 0 DDRB\[7\]
rlabel metal2 16408 43456 16408 43456 0 PORTA\[0\]
rlabel metal2 14728 39312 14728 39312 0 PORTA\[1\]
rlabel metal2 11088 43064 11088 43064 0 PORTA\[2\]
rlabel metal2 22344 42224 22344 42224 0 PORTA\[3\]
rlabel metal3 12936 38808 12936 38808 0 PORTA\[4\]
rlabel metal2 32368 39704 32368 39704 0 PORTA\[5\]
rlabel metal2 16856 40096 16856 40096 0 PORTA\[6\]
rlabel metal2 24584 34832 24584 34832 0 PORTA\[7\]
rlabel metal2 19656 30128 19656 30128 0 PORTB\[0\]
rlabel metal2 27608 32200 27608 32200 0 PORTB\[1\]
rlabel metal3 22232 26376 22232 26376 0 PORTB\[2\]
rlabel metal3 21000 34384 21000 34384 0 PORTB\[3\]
rlabel metal3 39928 37912 39928 37912 0 PORTB\[4\]
rlabel metal3 41440 34776 41440 34776 0 PORTB\[5\]
rlabel metal3 40320 42616 40320 42616 0 PORTB\[6\]
rlabel metal2 42616 31136 42616 31136 0 PORTB\[7\]
rlabel metal3 1358 35000 1358 35000 0 RXD
rlabel metal2 21448 36904 21448 36904 0 SPA\[0\]
rlabel metal2 14280 39312 14280 39312 0 SPA\[1\]
rlabel metal3 22680 34888 22680 34888 0 SPA\[2\]
rlabel metal2 27832 12712 27832 12712 0 SPA\[3\]
rlabel metal2 30016 12712 30016 12712 0 SPA\[4\]
rlabel metal2 29848 13720 29848 13720 0 SPA\[5\]
rlabel metal3 31024 12712 31024 12712 0 SPA\[6\]
rlabel metal2 10472 34944 10472 34944 0 SPA\[7\]
rlabel metal3 21728 26264 21728 26264 0 SPB\[0\]
rlabel metal2 31192 8036 31192 8036 0 SPB\[1\]
rlabel metal2 20440 25200 20440 25200 0 SPB\[2\]
rlabel metal3 29456 34776 29456 34776 0 SPB\[3\]
rlabel metal2 39256 15512 39256 15512 0 SPB\[4\]
rlabel metal3 39424 20216 39424 20216 0 SPB\[5\]
rlabel metal3 39704 19880 39704 19880 0 SPB\[6\]
rlabel metal2 41720 31248 41720 31248 0 SPB\[7\]
rlabel metal2 1736 33768 1736 33768 0 TXD
rlabel metal2 39816 27384 39816 27384 0 _000_
rlabel metal2 4480 21560 4480 21560 0 _001_
rlabel metal3 5712 22456 5712 22456 0 _002_
rlabel metal2 4984 25480 4984 25480 0 _003_
rlabel metal2 4312 27384 4312 27384 0 _004_
rlabel metal2 5096 28000 5096 28000 0 _005_
rlabel metal2 4256 28504 4256 28504 0 _006_
rlabel metal2 6104 31136 6104 31136 0 _007_
rlabel metal2 8008 31416 8008 31416 0 _008_
rlabel metal2 37800 24248 37800 24248 0 _009_
rlabel metal3 37464 26152 37464 26152 0 _010_
rlabel metal2 41272 24248 41272 24248 0 _011_
rlabel metal2 7336 38976 7336 38976 0 _012_
rlabel metal2 3080 36512 3080 36512 0 _013_
rlabel metal3 5992 41832 5992 41832 0 _014_
rlabel metal2 2744 40264 2744 40264 0 _015_
rlabel metal2 10584 42392 10584 42392 0 _016_
rlabel metal3 4928 36568 4928 36568 0 _017_
rlabel metal2 11816 42784 11816 42784 0 _018_
rlabel metal2 7392 44184 7392 44184 0 _019_
rlabel metal2 6776 15624 6776 15624 0 _020_
rlabel metal3 4872 17528 4872 17528 0 _021_
rlabel metal3 5488 16968 5488 16968 0 _022_
rlabel metal2 8232 12936 8232 12936 0 _023_
rlabel metal2 9464 10528 9464 10528 0 _024_
rlabel metal2 13384 9800 13384 9800 0 _025_
rlabel metal2 13720 11144 13720 11144 0 _026_
rlabel metal2 14840 14868 14840 14868 0 _027_
rlabel metal2 18088 11760 18088 11760 0 _028_
rlabel metal2 19544 8232 19544 8232 0 _029_
rlabel metal2 20888 6832 20888 6832 0 _030_
rlabel metal2 22568 14056 22568 14056 0 _031_
rlabel metal3 23184 8344 23184 8344 0 _032_
rlabel metal2 24248 13944 24248 13944 0 _033_
rlabel metal3 21672 16968 21672 16968 0 _034_
rlabel metal2 19376 17752 19376 17752 0 _035_
rlabel metal2 18424 43512 18424 43512 0 _036_
rlabel metal2 17752 42392 17752 42392 0 _037_
rlabel metal2 22568 43120 22568 43120 0 _038_
rlabel metal2 23464 42056 23464 42056 0 _039_
rlabel metal2 28056 41328 28056 41328 0 _040_
rlabel metal3 29176 39704 29176 39704 0 _041_
rlabel metal2 27608 39088 27608 39088 0 _042_
rlabel metal2 23912 38976 23912 38976 0 _043_
rlabel metal2 28336 29512 28336 29512 0 _044_
rlabel metal2 31864 30240 31864 30240 0 _045_
rlabel metal2 27496 27440 27496 27440 0 _046_
rlabel metal2 29288 33712 29288 33712 0 _047_
rlabel metal2 35560 34888 35560 34888 0 _048_
rlabel metal3 37240 33432 37240 33432 0 _049_
rlabel metal3 37296 32424 37296 32424 0 _050_
rlabel metal3 37744 30072 37744 30072 0 _051_
rlabel metal2 21896 31360 21896 31360 0 _052_
rlabel metal2 27944 18760 27944 18760 0 _053_
rlabel metal2 23352 26684 23352 26684 0 _054_
rlabel metal2 28504 11312 28504 11312 0 _055_
rlabel metal2 29960 10976 29960 10976 0 _056_
rlabel metal2 31752 11424 31752 11424 0 _057_
rlabel metal2 31304 13328 31304 13328 0 _058_
rlabel metal2 23744 30072 23744 30072 0 _059_
rlabel metal2 31136 23688 31136 23688 0 _060_
rlabel metal2 32760 16408 32760 16408 0 _061_
rlabel metal3 31640 20664 31640 20664 0 _062_
rlabel metal2 29736 24304 29736 24304 0 _063_
rlabel metal3 36456 15400 36456 15400 0 _064_
rlabel metal2 37800 16464 37800 16464 0 _065_
rlabel metal3 37240 19880 37240 19880 0 _066_
rlabel metal3 38248 20664 38248 20664 0 _067_
rlabel metal3 33208 35560 33208 35560 0 _068_
rlabel metal3 33208 27720 33208 27720 0 _069_
rlabel metal3 21000 43400 21000 43400 0 _070_
rlabel metal2 21000 43904 21000 43904 0 _071_
rlabel metal2 18816 39256 18816 39256 0 _072_
rlabel metal2 22064 17416 22064 17416 0 _073_
rlabel metal2 24360 44016 24360 44016 0 _074_
rlabel metal2 28896 37464 28896 37464 0 _075_
rlabel metal2 30408 40096 30408 40096 0 _076_
rlabel metal3 32984 40264 32984 40264 0 _077_
rlabel metal2 34048 39032 34048 39032 0 _078_
rlabel metal3 19824 25928 19824 25928 0 _079_
rlabel metal3 31640 41384 31640 41384 0 _080_
rlabel metal2 17976 24808 17976 24808 0 _081_
rlabel metal2 20496 23240 20496 23240 0 _082_
rlabel metal3 35280 43512 35280 43512 0 _083_
rlabel metal2 35672 41496 35672 41496 0 _084_
rlabel metal3 23968 6664 23968 6664 0 _085_
rlabel metal2 26264 27160 26264 27160 0 _086_
rlabel metal2 25592 23520 25592 23520 0 _087_
rlabel metal3 32032 44184 32032 44184 0 _088_
rlabel metal2 40152 38416 40152 38416 0 _089_
rlabel metal2 41608 35784 41608 35784 0 _090_
rlabel metal3 42392 44184 42392 44184 0 _091_
rlabel metal2 43512 37688 43512 37688 0 _092_
rlabel metal2 19208 24192 19208 24192 0 _093_
rlabel metal2 22568 5320 22568 5320 0 _094_
rlabel metal3 30464 43512 30464 43512 0 _095_
rlabel metal2 44632 43120 44632 43120 0 _096_
rlabel metal2 10808 28280 10808 28280 0 _097_
rlabel metal3 11144 38808 11144 38808 0 _098_
rlabel metal2 39704 24752 39704 24752 0 _099_
rlabel metal2 38808 28392 38808 28392 0 _100_
rlabel metal2 19880 21616 19880 21616 0 _101_
rlabel metal3 11984 32536 11984 32536 0 _102_
rlabel metal2 9912 31920 9912 31920 0 _103_
rlabel metal2 7224 24864 7224 24864 0 _104_
rlabel metal2 5992 23072 5992 23072 0 _105_
rlabel metal3 11312 19880 11312 19880 0 _106_
rlabel metal2 15568 18536 15568 18536 0 _107_
rlabel metal3 13048 19208 13048 19208 0 _108_
rlabel metal2 12544 19432 12544 19432 0 _109_
rlabel metal2 18032 23352 18032 23352 0 _110_
rlabel metal2 19768 30576 19768 30576 0 _111_
rlabel metal2 12600 21448 12600 21448 0 _112_
rlabel metal2 12712 23072 12712 23072 0 _113_
rlabel metal2 11704 22736 11704 22736 0 _114_
rlabel metal2 18088 23128 18088 23128 0 _115_
rlabel metal2 12824 19768 12824 19768 0 _116_
rlabel metal2 15400 21392 15400 21392 0 _117_
rlabel metal3 15204 23240 15204 23240 0 _118_
rlabel metal2 15176 25200 15176 25200 0 _119_
rlabel metal2 21224 26208 21224 26208 0 _120_
rlabel metal3 12320 24696 12320 24696 0 _121_
rlabel metal2 13776 32536 13776 32536 0 _122_
rlabel metal3 18368 26488 18368 26488 0 _123_
rlabel metal3 19880 26152 19880 26152 0 _124_
rlabel metal2 13440 24808 13440 24808 0 _125_
rlabel metal2 21560 21280 21560 21280 0 _126_
rlabel metal3 24248 23800 24248 23800 0 _127_
rlabel metal2 18984 32200 18984 32200 0 _128_
rlabel metal3 17752 29400 17752 29400 0 _129_
rlabel metal2 17416 23408 17416 23408 0 _130_
rlabel metal3 9912 21560 9912 21560 0 _131_
rlabel metal2 10080 22456 10080 22456 0 _132_
rlabel metal3 13328 38696 13328 38696 0 _133_
rlabel metal2 16408 22792 16408 22792 0 _134_
rlabel metal2 16632 23296 16632 23296 0 _135_
rlabel metal2 14616 39200 14616 39200 0 _136_
rlabel metal2 24808 21112 24808 21112 0 _137_
rlabel metal2 16744 39144 16744 39144 0 _138_
rlabel metal2 15400 32816 15400 32816 0 _139_
rlabel metal3 15400 39704 15400 39704 0 _140_
rlabel metal2 15624 21056 15624 21056 0 _141_
rlabel metal2 15176 19768 15176 19768 0 _142_
rlabel metal2 9016 23576 9016 23576 0 _143_
rlabel metal2 19040 34104 19040 34104 0 _144_
rlabel metal3 14616 31136 14616 31136 0 _145_
rlabel metal2 8232 24360 8232 24360 0 _146_
rlabel metal2 8624 23688 8624 23688 0 _147_
rlabel metal3 6608 23128 6608 23128 0 _148_
rlabel metal2 12376 32592 12376 32592 0 _149_
rlabel metal2 9016 22120 9016 22120 0 _150_
rlabel metal2 7784 23072 7784 23072 0 _151_
rlabel metal2 14280 35224 14280 35224 0 _152_
rlabel metal2 14056 34664 14056 34664 0 _153_
rlabel metal2 19432 31304 19432 31304 0 _154_
rlabel metal2 19432 25480 19432 25480 0 _155_
rlabel metal2 13944 32984 13944 32984 0 _156_
rlabel metal2 3192 29120 3192 29120 0 _157_
rlabel metal3 7560 25704 7560 25704 0 _158_
rlabel metal2 18424 22176 18424 22176 0 _159_
rlabel metal2 18312 24360 18312 24360 0 _160_
rlabel metal2 18536 25032 18536 25032 0 _161_
rlabel metal2 8680 25760 8680 25760 0 _162_
rlabel metal2 16408 36008 16408 36008 0 _163_
rlabel metal2 10248 37520 10248 37520 0 _164_
rlabel metal2 10024 36904 10024 36904 0 _165_
rlabel metal2 9128 31976 9128 31976 0 _166_
rlabel metal2 13552 38696 13552 38696 0 _167_
rlabel metal2 8904 31640 8904 31640 0 _168_
rlabel metal2 8904 27104 8904 27104 0 _169_
rlabel metal2 8512 27608 8512 27608 0 _170_
rlabel metal2 9464 30520 9464 30520 0 _171_
rlabel metal3 7616 27272 7616 27272 0 _172_
rlabel metal3 18144 27944 18144 27944 0 _173_
rlabel metal2 17528 27160 17528 27160 0 _174_
rlabel metal3 16044 26824 16044 26824 0 _175_
rlabel metal2 15960 35728 15960 35728 0 _176_
rlabel metal3 11032 34776 11032 34776 0 _177_
rlabel metal2 8848 34888 8848 34888 0 _178_
rlabel metal2 9016 28224 9016 28224 0 _179_
rlabel metal3 8792 27720 8792 27720 0 _180_
rlabel metal2 17192 24472 17192 24472 0 _181_
rlabel metal3 1848 44296 1848 44296 0 _182_
rlabel metal2 16632 25312 16632 25312 0 _183_
rlabel metal3 12320 26824 12320 26824 0 _184_
rlabel metal2 12040 38136 12040 38136 0 _185_
rlabel metal2 19208 36120 19208 36120 0 _186_
rlabel metal2 10416 27944 10416 27944 0 _187_
rlabel metal3 8400 28616 8400 28616 0 _188_
rlabel metal2 18200 28448 18200 28448 0 _189_
rlabel metal2 12040 32928 12040 32928 0 _190_
rlabel metal3 12768 35336 12768 35336 0 _191_
rlabel metal2 11704 35448 11704 35448 0 _192_
rlabel metal2 12040 33768 12040 33768 0 _193_
rlabel metal2 9912 29904 9912 29904 0 _194_
rlabel metal3 8792 30968 8792 30968 0 _195_
rlabel metal2 10248 30632 10248 30632 0 _196_
rlabel metal2 16800 38696 16800 38696 0 _197_
rlabel metal2 18200 33488 18200 33488 0 _198_
rlabel metal2 19208 31472 19208 31472 0 _199_
rlabel metal2 10584 31640 10584 31640 0 _200_
rlabel metal2 8120 31304 8120 31304 0 _201_
rlabel metal2 1512 36848 1512 36848 0 _202_
rlabel metal3 13888 26488 13888 26488 0 _203_
rlabel metal2 15176 29792 15176 29792 0 _204_
rlabel metal3 11704 29960 11704 29960 0 _205_
rlabel metal2 9632 35448 9632 35448 0 _206_
rlabel metal3 13496 25592 13496 25592 0 _207_
rlabel metal2 11928 31304 11928 31304 0 _208_
rlabel metal2 9128 31024 9128 31024 0 _209_
rlabel metal2 21784 22848 21784 22848 0 _210_
rlabel metal3 22904 21560 22904 21560 0 _211_
rlabel metal3 22288 21672 22288 21672 0 _212_
rlabel metal2 23464 23968 23464 23968 0 _213_
rlabel metal2 34664 25704 34664 25704 0 _214_
rlabel metal2 32200 36008 32200 36008 0 _215_
rlabel metal2 35448 25480 35448 25480 0 _216_
rlabel metal2 36344 25088 36344 25088 0 _217_
rlabel metal2 34440 25928 34440 25928 0 _218_
rlabel metal3 35224 26712 35224 26712 0 _219_
rlabel metal2 32200 28224 32200 28224 0 _220_
rlabel metal2 35224 27048 35224 27048 0 _221_
rlabel metal2 36344 26264 36344 26264 0 _222_
rlabel metal2 23800 20384 23800 20384 0 _223_
rlabel metal2 35000 25200 35000 25200 0 _224_
rlabel metal2 39592 25984 39592 25984 0 _225_
rlabel metal2 39480 24752 39480 24752 0 _226_
rlabel metal2 9016 40656 9016 40656 0 _227_
rlabel metal2 15736 23912 15736 23912 0 _228_
rlabel metal2 18704 22456 18704 22456 0 _229_
rlabel metal3 13664 40376 13664 40376 0 _230_
rlabel metal2 8568 40768 8568 40768 0 _231_
rlabel metal2 7168 39592 7168 39592 0 _232_
rlabel metal2 23912 23016 23912 23016 0 _233_
rlabel metal2 8176 39144 8176 39144 0 _234_
rlabel metal2 4144 34216 4144 34216 0 _235_
rlabel metal3 3332 38024 3332 38024 0 _236_
rlabel metal3 6048 39480 6048 39480 0 _237_
rlabel metal2 7336 40040 7336 40040 0 _238_
rlabel metal2 3864 35560 3864 35560 0 _239_
rlabel metal3 3248 34888 3248 34888 0 _240_
rlabel metal2 3304 34720 3304 34720 0 _241_
rlabel metal3 10976 41272 10976 41272 0 _242_
rlabel metal3 8008 41944 8008 41944 0 _243_
rlabel metal2 8120 41720 8120 41720 0 _244_
rlabel metal2 7672 42224 7672 42224 0 _245_
rlabel metal2 4984 37128 4984 37128 0 _246_
rlabel metal2 3752 36008 3752 36008 0 _247_
rlabel metal2 12488 14504 12488 14504 0 _248_
rlabel metal3 11368 41384 11368 41384 0 _249_
rlabel metal2 10248 42000 10248 42000 0 _250_
rlabel metal2 2968 37240 2968 37240 0 _251_
rlabel metal2 4816 35112 4816 35112 0 _252_
rlabel metal2 24360 21840 24360 21840 0 _253_
rlabel metal2 23800 22568 23800 22568 0 _254_
rlabel metal2 13720 40768 13720 40768 0 _255_
rlabel metal2 12488 41440 12488 41440 0 _256_
rlabel metal2 10640 43288 10640 43288 0 _257_
rlabel metal2 14392 40712 14392 40712 0 _258_
rlabel metal2 8232 41888 8232 41888 0 _259_
rlabel metal2 7896 42784 7896 42784 0 _260_
rlabel metal2 11256 14224 11256 14224 0 _261_
rlabel metal3 8904 42056 8904 42056 0 _262_
rlabel metal3 20664 21784 20664 21784 0 _263_
rlabel metal2 15736 18144 15736 18144 0 _264_
rlabel metal2 10696 16184 10696 16184 0 _265_
rlabel metal3 7448 16072 7448 16072 0 _266_
rlabel metal3 13888 15512 13888 15512 0 _267_
rlabel metal2 6104 16800 6104 16800 0 _268_
rlabel metal2 6552 15960 6552 15960 0 _269_
rlabel metal2 19320 40656 19320 40656 0 _270_
rlabel metal3 7728 17528 7728 17528 0 _271_
rlabel metal2 6552 17528 6552 17528 0 _272_
rlabel metal3 8064 16968 8064 16968 0 _273_
rlabel metal2 7560 17024 7560 17024 0 _274_
rlabel metal2 26544 15176 26544 15176 0 _275_
rlabel metal2 9968 13832 9968 13832 0 _276_
rlabel metal2 9632 13832 9632 13832 0 _277_
rlabel metal2 13944 12600 13944 12600 0 _278_
rlabel metal2 14336 14504 14336 14504 0 _279_
rlabel metal2 11704 13272 11704 13272 0 _280_
rlabel metal2 12712 13384 12712 13384 0 _281_
rlabel metal2 11928 12600 11928 12600 0 _282_
rlabel metal2 14392 14280 14392 14280 0 _283_
rlabel metal2 13720 12264 13720 12264 0 _284_
rlabel metal2 14112 12152 14112 12152 0 _285_
rlabel metal2 13720 13048 13720 13048 0 _286_
rlabel metal2 13216 12936 13216 12936 0 _287_
rlabel metal2 15064 15176 15064 15176 0 _288_
rlabel metal2 15624 15624 15624 15624 0 _289_
rlabel metal3 21784 14504 21784 14504 0 _290_
rlabel metal2 18200 18648 18200 18648 0 _291_
rlabel metal2 21448 16408 21448 16408 0 _292_
rlabel metal2 18984 12768 18984 12768 0 _293_
rlabel metal2 20664 15680 20664 15680 0 _294_
rlabel metal2 21672 11928 21672 11928 0 _295_
rlabel metal2 21896 10248 21896 10248 0 _296_
rlabel metal2 19264 10808 19264 10808 0 _297_
rlabel metal2 19544 9184 19544 9184 0 _298_
rlabel metal2 19320 9464 19320 9464 0 _299_
rlabel metal2 20944 9016 20944 9016 0 _300_
rlabel metal2 19880 14896 19880 14896 0 _301_
rlabel metal2 19712 16968 19712 16968 0 _302_
rlabel metal2 21224 14280 21224 14280 0 _303_
rlabel metal2 22344 10752 22344 10752 0 _304_
rlabel metal3 21896 15288 21896 15288 0 _305_
rlabel metal3 20496 15288 20496 15288 0 _306_
rlabel metal2 21056 16856 21056 16856 0 _307_
rlabel metal3 20216 16968 20216 16968 0 _308_
rlabel metal2 17080 21112 17080 21112 0 _309_
rlabel metal2 19544 17920 19544 17920 0 _310_
rlabel metal2 19208 18312 19208 18312 0 _311_
rlabel metal3 20496 39368 20496 39368 0 _312_
rlabel metal3 22848 41048 22848 41048 0 _313_
rlabel metal2 18648 42000 18648 42000 0 _314_
rlabel metal2 20328 40040 20328 40040 0 _315_
rlabel via2 18536 42168 18536 42168 0 _316_
rlabel metal2 18200 42672 18200 42672 0 _317_
rlabel metal2 17808 41160 17808 41160 0 _318_
rlabel metal2 18200 42000 18200 42000 0 _319_
rlabel metal2 23296 41384 23296 41384 0 _320_
rlabel metal2 22232 42728 22232 42728 0 _321_
rlabel metal3 29064 39032 29064 39032 0 _322_
rlabel metal2 23912 41888 23912 41888 0 _323_
rlabel metal2 22904 41272 22904 41272 0 _324_
rlabel metal2 22680 41944 22680 41944 0 _325_
rlabel metal3 22064 39368 22064 39368 0 _326_
rlabel metal2 27832 40824 27832 40824 0 _327_
rlabel metal2 22344 39536 22344 39536 0 _328_
rlabel metal2 28392 40880 28392 40880 0 _329_
rlabel metal2 27272 38976 27272 38976 0 _330_
rlabel metal2 27776 39592 27776 39592 0 _331_
rlabel metal2 27720 38640 27720 38640 0 _332_
rlabel metal2 27496 39256 27496 39256 0 _333_
rlabel metal2 24024 39200 24024 39200 0 _334_
rlabel metal3 23296 39480 23296 39480 0 _335_
rlabel metal2 23352 38920 23352 38920 0 _336_
rlabel metal2 25592 30912 25592 30912 0 _337_
rlabel metal2 29064 31808 29064 31808 0 _338_
rlabel metal3 28392 30968 28392 30968 0 _339_
rlabel metal3 24472 25816 24472 25816 0 _340_
rlabel metal2 26488 27832 26488 27832 0 _341_
rlabel metal2 27664 31080 27664 31080 0 _342_
rlabel metal2 27048 32368 27048 32368 0 _343_
rlabel metal2 27944 32536 27944 32536 0 _344_
rlabel metal2 25928 27160 25928 27160 0 _345_
rlabel metal2 23800 26264 23800 26264 0 _346_
rlabel metal3 28560 33320 28560 33320 0 _347_
rlabel metal2 29064 33264 29064 33264 0 _348_
rlabel metal3 30072 33208 30072 33208 0 _349_
rlabel metal2 29456 32760 29456 32760 0 _350_
rlabel metal2 34776 32256 34776 32256 0 _351_
rlabel metal2 35000 33824 35000 33824 0 _352_
rlabel metal2 34104 30744 34104 30744 0 _353_
rlabel metal2 35112 33040 35112 33040 0 _354_
rlabel metal2 36176 31192 36176 31192 0 _355_
rlabel metal2 35672 32592 35672 32592 0 _356_
rlabel metal2 35224 29680 35224 29680 0 _357_
rlabel metal2 36008 30464 36008 30464 0 _358_
rlabel metal3 27664 12152 27664 12152 0 _359_
rlabel metal2 25032 21448 25032 21448 0 _360_
rlabel metal2 23800 24640 23800 24640 0 _361_
rlabel metal3 25200 24808 25200 24808 0 _362_
rlabel metal3 22736 27272 22736 27272 0 _363_
rlabel metal2 26040 18592 26040 18592 0 _364_
rlabel metal2 28056 14056 28056 14056 0 _365_
rlabel metal2 27272 18368 27272 18368 0 _366_
rlabel metal2 26768 19208 26768 19208 0 _367_
rlabel metal2 24136 26096 24136 26096 0 _368_
rlabel metal2 27664 12152 27664 12152 0 _369_
rlabel metal2 27832 13160 27832 13160 0 _370_
rlabel metal2 27496 12488 27496 12488 0 _371_
rlabel metal2 29624 12432 29624 12432 0 _372_
rlabel metal2 29792 12264 29792 12264 0 _373_
rlabel metal2 30520 14504 30520 14504 0 _374_
rlabel metal2 30184 13832 30184 13832 0 _375_
rlabel metal3 31248 13832 31248 13832 0 _376_
rlabel metal2 31416 14420 31416 14420 0 _377_
rlabel metal2 30856 12936 30856 12936 0 _378_
rlabel metal3 23744 27048 23744 27048 0 _379_
rlabel metal2 29624 22232 29624 22232 0 _380_
rlabel metal2 30128 23800 30128 23800 0 _381_
rlabel metal2 30520 23016 30520 23016 0 _382_
rlabel metal2 25928 20216 25928 20216 0 _383_
rlabel metal2 31752 19432 31752 19432 0 _384_
rlabel metal2 31192 17136 31192 17136 0 _385_
rlabel metal2 31248 17640 31248 17640 0 _386_
rlabel metal2 30464 20216 30464 20216 0 _387_
rlabel metal3 29680 20776 29680 20776 0 _388_
rlabel metal2 27608 23632 27608 23632 0 _389_
rlabel metal2 31752 16520 31752 16520 0 _390_
rlabel metal3 35560 19208 35560 19208 0 _391_
rlabel metal2 36008 16576 36008 16576 0 _392_
rlabel metal2 36680 16968 36680 16968 0 _393_
rlabel metal3 34944 16856 34944 16856 0 _394_
rlabel metal2 36288 16968 36288 16968 0 _395_
rlabel metal3 35896 19992 35896 19992 0 _396_
rlabel metal2 36344 19712 36344 19712 0 _397_
rlabel metal2 35784 20160 35784 20160 0 _398_
rlabel metal2 37128 20272 37128 20272 0 _399_
rlabel metal2 1736 2744 1736 2744 0 addr[0]
rlabel metal2 1736 3976 1736 3976 0 addr[1]
rlabel metal3 1302 5208 1302 5208 0 addr[2]
rlabel metal2 1736 7112 1736 7112 0 addr[3]
rlabel metal2 35392 3416 35392 3416 0 bus_cyc
rlabel metal2 37016 2086 37016 2086 0 bus_we
rlabel metal2 28952 14224 28952 14224 0 clknet_0_wb_clk_i
rlabel metal2 14840 9408 14840 9408 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 2520 16072 2520 16072 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 29176 11144 29176 11144 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 40152 23632 40152 23632 0 clknet_3_3__leaf_wb_clk_i
rlabel metal2 8120 38920 8120 38920 0 clknet_3_4__leaf_wb_clk_i
rlabel metal3 5432 44296 5432 44296 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 38920 30072 38920 30072 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 25368 42728 25368 42728 0 clknet_3_7__leaf_wb_clk_i
rlabel metal3 1246 8344 1246 8344 0 data_in[0]
rlabel metal3 1302 9912 1302 9912 0 data_in[1]
rlabel metal3 1302 11480 1302 11480 0 data_in[2]
rlabel metal3 1302 13048 1302 13048 0 data_in[3]
rlabel metal2 1736 14560 1736 14560 0 data_in[4]
rlabel metal3 1302 16184 1302 16184 0 data_in[5]
rlabel metal2 1736 18088 1736 18088 0 data_in[6]
rlabel metal2 1736 19656 1736 19656 0 data_in[7]
rlabel metal3 1358 20888 1358 20888 0 data_out[0]
rlabel metal3 1358 22456 1358 22456 0 data_out[1]
rlabel metal3 1358 24024 1358 24024 0 data_out[2]
rlabel metal3 1358 25592 1358 25592 0 data_out[3]
rlabel metal3 1358 27160 1358 27160 0 data_out[4]
rlabel metal3 1358 28728 1358 28728 0 data_out[5]
rlabel metal3 1358 30296 1358 30296 0 data_out[6]
rlabel metal3 1302 31864 1302 31864 0 data_out[7]
rlabel metal2 5656 46368 5656 46368 0 io_in[0]
rlabel metal2 16296 45976 16296 45976 0 io_in[10]
rlabel metal2 17640 45864 17640 45864 0 io_in[11]
rlabel metal2 18872 47642 18872 47642 0 io_in[12]
rlabel metal2 20216 47642 20216 47642 0 io_in[13]
rlabel metal2 22008 45976 22008 45976 0 io_in[14]
rlabel metal2 22904 47642 22904 47642 0 io_in[15]
rlabel metal2 4424 44408 4424 44408 0 io_in[1]
rlabel metal3 5096 45864 5096 45864 0 io_in[2]
rlabel metal2 7224 46368 7224 46368 0 io_in[3]
rlabel metal2 8120 47642 8120 47642 0 io_in[4]
rlabel metal2 9576 45864 9576 45864 0 io_in[5]
rlabel metal2 10808 47642 10808 47642 0 io_in[6]
rlabel metal2 12208 45864 12208 45864 0 io_in[7]
rlabel metal2 13496 47642 13496 47642 0 io_in[8]
rlabel metal2 14840 47642 14840 47642 0 io_in[9]
rlabel metal2 2744 2198 2744 2198 0 io_oeb[0]
rlabel metal2 22904 1582 22904 1582 0 io_oeb[10]
rlabel metal2 24920 2058 24920 2058 0 io_oeb[11]
rlabel metal2 26936 2422 26936 2422 0 io_oeb[12]
rlabel metal2 28952 2086 28952 2086 0 io_oeb[13]
rlabel metal2 30968 2086 30968 2086 0 io_oeb[14]
rlabel metal2 32984 2422 32984 2422 0 io_oeb[15]
rlabel metal2 4760 2030 4760 2030 0 io_oeb[1]
rlabel metal2 6776 2198 6776 2198 0 io_oeb[2]
rlabel metal2 8792 2422 8792 2422 0 io_oeb[3]
rlabel metal2 10808 2086 10808 2086 0 io_oeb[4]
rlabel metal2 12824 2422 12824 2422 0 io_oeb[5]
rlabel metal2 14840 2086 14840 2086 0 io_oeb[6]
rlabel metal2 16856 854 16856 854 0 io_oeb[7]
rlabel metal2 18872 2058 18872 2058 0 io_oeb[8]
rlabel metal3 21504 3640 21504 3640 0 io_oeb[9]
rlabel metal2 24248 46914 24248 46914 0 io_out[0]
rlabel metal2 37688 47698 37688 47698 0 io_out[10]
rlabel metal2 39032 46914 39032 46914 0 io_out[11]
rlabel metal2 40376 47306 40376 47306 0 io_out[12]
rlabel metal2 41720 47698 41720 47698 0 io_out[13]
rlabel metal2 43064 47306 43064 47306 0 io_out[14]
rlabel metal2 44408 46914 44408 46914 0 io_out[15]
rlabel metal2 26264 47712 26264 47712 0 io_out[1]
rlabel metal2 26936 47306 26936 47306 0 io_out[2]
rlabel metal2 28280 47698 28280 47698 0 io_out[3]
rlabel metal2 29624 46914 29624 46914 0 io_out[4]
rlabel metal2 30968 47698 30968 47698 0 io_out[5]
rlabel metal2 32312 47138 32312 47138 0 io_out[6]
rlabel metal2 33656 47698 33656 47698 0 io_out[7]
rlabel metal2 35000 47306 35000 47306 0 io_out[8]
rlabel metal3 37184 44520 37184 44520 0 io_out[9]
rlabel metal2 39032 2198 39032 2198 0 irq0
rlabel metal2 41048 2422 41048 2422 0 irq6
rlabel metal2 43064 854 43064 854 0 irq7
rlabel metal3 1358 36568 1358 36568 0 la_data_out[0]
rlabel metal3 1358 38136 1358 38136 0 la_data_out[1]
rlabel metal3 1358 39704 1358 39704 0 la_data_out[2]
rlabel metal3 1414 41272 1414 41272 0 la_data_out[3]
rlabel metal3 1358 42840 1358 42840 0 la_data_out[4]
rlabel metal3 1302 44408 1302 44408 0 la_data_out[5]
rlabel metal3 1358 45976 1358 45976 0 la_data_out[6]
rlabel metal3 2814 47544 2814 47544 0 la_data_out[7]
rlabel metal3 35504 27720 35504 27720 0 last_irg6_trigger
rlabel metal2 35112 35224 35112 35224 0 last_irq0_trigger
rlabel metal2 41944 27496 41944 27496 0 last_irq7_trigger
rlabel metal2 43176 31024 43176 31024 0 net1
rlabel metal2 36008 4200 36008 4200 0 net10
rlabel metal2 4312 40320 4312 40320 0 net100
rlabel metal2 7224 45360 7224 45360 0 net101
rlabel metal3 5264 44072 5264 44072 0 net102
rlabel metal3 5880 42616 5880 42616 0 net103
rlabel metal2 23352 18144 23352 18144 0 net11
rlabel metal3 3808 9240 3808 9240 0 net12
rlabel metal3 2688 10696 2688 10696 0 net13
rlabel metal3 5348 12040 5348 12040 0 net14
rlabel metal3 2912 13720 2912 13720 0 net15
rlabel metal2 2408 12992 2408 12992 0 net16
rlabel metal2 2296 17136 2296 17136 0 net17
rlabel metal2 2072 18368 2072 18368 0 net18
rlabel metal2 2072 19936 2072 19936 0 net19
rlabel metal3 47880 36120 47880 36120 0 net2
rlabel metal2 19544 26488 19544 26488 0 net20
rlabel metal2 17304 44240 17304 44240 0 net21
rlabel metal3 19096 43288 19096 43288 0 net22
rlabel metal3 18704 45416 18704 45416 0 net23
rlabel metal3 20104 41944 20104 41944 0 net24
rlabel metal3 20384 45752 20384 45752 0 net25
rlabel metal2 15288 45024 15288 45024 0 net26
rlabel metal2 11592 36624 11592 36624 0 net27
rlabel metal3 6216 43960 6216 43960 0 net28
rlabel metal3 8148 45192 8148 45192 0 net29
rlabel metal2 47880 39480 47880 39480 0 net3
rlabel metal2 14728 44744 14728 44744 0 net30
rlabel metal2 9912 45640 9912 45640 0 net31
rlabel metal2 11312 45640 11312 45640 0 net32
rlabel metal2 12600 44660 12600 44660 0 net33
rlabel metal2 17416 30240 17416 30240 0 net34
rlabel metal2 15400 42672 15400 42672 0 net35
rlabel metal3 41888 14280 41888 14280 0 net36
rlabel metal3 47040 20104 47040 20104 0 net37
rlabel metal2 47880 25424 47880 25424 0 net38
rlabel metal3 47096 3640 47096 3640 0 net39
rlabel metal2 47880 45024 47880 45024 0 net4
rlabel metal3 46200 4536 46200 4536 0 net40
rlabel metal3 40096 9128 40096 9128 0 net41
rlabel metal3 5824 35112 5824 35112 0 net42
rlabel metal2 2296 21112 2296 21112 0 net43
rlabel metal2 2072 22792 2072 22792 0 net44
rlabel metal3 5544 23912 5544 23912 0 net45
rlabel metal2 2184 27048 2184 27048 0 net46
rlabel metal2 2968 27664 2968 27664 0 net47
rlabel metal2 4312 29064 4312 29064 0 net48
rlabel metal3 5824 30856 5824 30856 0 net49
rlabel metal2 2072 34888 2072 34888 0 net5
rlabel metal2 1960 31808 1960 31808 0 net50
rlabel metal2 5208 11816 5208 11816 0 net51
rlabel metal2 22792 5040 22792 5040 0 net52
rlabel metal3 27888 3528 27888 3528 0 net53
rlabel metal2 27160 6356 27160 6356 0 net54
rlabel metal3 28672 5992 28672 5992 0 net55
rlabel metal3 33152 3528 33152 3528 0 net56
rlabel metal2 33208 6356 33208 6356 0 net57
rlabel metal3 6552 15960 6552 15960 0 net58
rlabel metal2 8232 17752 8232 17752 0 net59
rlabel metal2 2016 3416 2016 3416 0 net6
rlabel metal2 12040 7336 12040 7336 0 net60
rlabel metal2 12600 6552 12600 6552 0 net61
rlabel metal2 13384 6356 13384 6356 0 net62
rlabel metal2 16016 11256 16016 11256 0 net63
rlabel metal3 18536 3528 18536 3528 0 net64
rlabel metal2 21672 6720 21672 6720 0 net65
rlabel metal2 21336 5376 21336 5376 0 net66
rlabel metal2 22792 44240 22792 44240 0 net67
rlabel metal2 39816 45696 39816 45696 0 net68
rlabel metal2 39928 44240 39928 44240 0 net69
rlabel metal2 2072 5096 2072 5096 0 net7
rlabel metal2 39816 40432 39816 40432 0 net70
rlabel metal2 43960 41048 43960 41048 0 net71
rlabel metal2 43176 44632 43176 44632 0 net72
rlabel metal2 43848 44240 43848 44240 0 net73
rlabel metal2 24136 45024 24136 45024 0 net74
rlabel metal3 26404 45192 26404 45192 0 net75
rlabel metal2 29176 45024 29176 45024 0 net76
rlabel metal2 29960 44016 29960 44016 0 net77
rlabel metal2 31864 45584 31864 45584 0 net78
rlabel metal2 34440 44632 34440 44632 0 net79
rlabel metal2 2464 5880 2464 5880 0 net8
rlabel metal2 33096 45024 33096 45024 0 net80
rlabel metal2 33432 43680 33432 43680 0 net81
rlabel metal2 35672 44240 35672 44240 0 net82
rlabel metal2 42056 4256 42056 4256 0 net83
rlabel metal2 40320 4536 40320 4536 0 net84
rlabel metal3 46200 3528 46200 3528 0 net85
rlabel metal2 5152 38696 5152 38696 0 net86
rlabel metal2 8064 37240 8064 37240 0 net87
rlabel metal2 6664 41160 6664 41160 0 net88
rlabel metal3 5208 41272 5208 41272 0 net89
rlabel metal2 2072 8036 2072 8036 0 net9
rlabel metal2 11704 43876 11704 43876 0 net90
rlabel metal2 1960 44044 1960 44044 0 net91
rlabel metal2 14280 41496 14280 41496 0 net92
rlabel metal2 8120 43232 8120 43232 0 net93
rlabel metal3 42140 43512 42140 43512 0 net94
rlabel metal2 45304 43176 45304 43176 0 net95
rlabel metal2 4312 45696 4312 45696 0 net96
rlabel metal2 7672 37744 7672 37744 0 net97
rlabel metal3 5544 42728 5544 42728 0 net98
rlabel metal2 4312 36792 4312 36792 0 net99
rlabel metal2 48216 14280 48216 14280 0 pwm0
rlabel metal2 48216 19768 48216 19768 0 pwm1
rlabel metal2 48216 25144 48216 25144 0 pwm2
rlabel metal2 47432 2968 47432 2968 0 rst
rlabel metal3 46200 43400 46200 43400 0 tmr0_clk
rlabel metal2 48216 3864 48216 3864 0 tmr0_o
rlabel metal2 47096 46130 47096 46130 0 tmr1_clk
rlabel metal2 48216 8904 48216 8904 0 tmr1_o
rlabel metal2 45080 13006 45080 13006 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
