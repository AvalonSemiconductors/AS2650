// This is the unpowered netlist.
module wrapped_as2650 (WEb_raw,
    boot_rom_en,
    bus_cyc,
    bus_we_gpios,
    bus_we_serial_ports,
    bus_we_sid,
    bus_we_timers,
    le_hi_act,
    le_lo_act,
    ram_enabled,
    reset_out,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    RAM_end_addr,
    RAM_start_addr,
    bus_addr,
    bus_data_out,
    bus_in_gpios,
    bus_in_serial_ports,
    bus_in_sid,
    bus_in_timers,
    cs_port,
    io_in,
    io_oeb,
    io_out,
    irq,
    irqs,
    la_data_out,
    last_addr,
    ram_bus_in,
    requested_addr,
    rom_bus_in,
    rom_bus_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output WEb_raw;
 output boot_rom_en;
 output bus_cyc;
 output bus_we_gpios;
 output bus_we_serial_ports;
 output bus_we_sid;
 output bus_we_timers;
 output le_hi_act;
 output le_lo_act;
 output ram_enabled;
 output reset_out;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [15:0] RAM_end_addr;
 output [15:0] RAM_start_addr;
 output [5:0] bus_addr;
 output [7:0] bus_data_out;
 input [7:0] bus_in_gpios;
 input [7:0] bus_in_serial_ports;
 input [7:0] bus_in_sid;
 input [7:0] bus_in_timers;
 output [2:0] cs_port;
 input [18:0] io_in;
 output [18:0] io_oeb;
 output [18:0] io_out;
 output [2:0] irq;
 input [6:0] irqs;
 output [55:0] la_data_out;
 output [15:0] last_addr;
 input [7:0] ram_bus_in;
 output [15:0] requested_addr;
 input [7:0] rom_bus_in;
 output [7:0] rom_bus_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire net331;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net310;
 wire net311;
 wire net332;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire \as2650.PC[0] ;
 wire \as2650.PC[10] ;
 wire \as2650.PC[11] ;
 wire \as2650.PC[12] ;
 wire \as2650.PC[1] ;
 wire \as2650.PC[2] ;
 wire \as2650.PC[3] ;
 wire \as2650.PC[4] ;
 wire \as2650.PC[5] ;
 wire \as2650.PC[6] ;
 wire \as2650.PC[7] ;
 wire \as2650.PC[8] ;
 wire \as2650.PC[9] ;
 wire \as2650.chirp_ptr[0] ;
 wire \as2650.chirp_ptr[1] ;
 wire \as2650.chirp_ptr[2] ;
 wire \as2650.chirpchar[0] ;
 wire \as2650.chirpchar[1] ;
 wire \as2650.chirpchar[2] ;
 wire \as2650.chirpchar[3] ;
 wire \as2650.chirpchar[4] ;
 wire \as2650.chirpchar[5] ;
 wire \as2650.chirpchar[6] ;
 wire \as2650.cpu_hidden_rom_enable ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[10] ;
 wire \as2650.cycle[11] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.cycle[8] ;
 wire \as2650.cycle[9] ;
 wire \as2650.debug_psl[0] ;
 wire \as2650.debug_psl[1] ;
 wire \as2650.debug_psl[2] ;
 wire \as2650.debug_psl[3] ;
 wire \as2650.debug_psl[4] ;
 wire \as2650.debug_psl[5] ;
 wire \as2650.debug_psl[6] ;
 wire \as2650.debug_psl[7] ;
 wire \as2650.debug_psu[0] ;
 wire \as2650.debug_psu[1] ;
 wire \as2650.debug_psu[2] ;
 wire \as2650.debug_psu[3] ;
 wire \as2650.debug_psu[4] ;
 wire \as2650.debug_psu[5] ;
 wire \as2650.debug_psu[7] ;
 wire \as2650.ext_io_addr[6] ;
 wire \as2650.ext_io_addr[7] ;
 wire \as2650.extend ;
 wire \as2650.indexed_cyc[0] ;
 wire \as2650.indexed_cyc[1] ;
 wire \as2650.indirect_cyc ;
 wire \as2650.indirect_target[0] ;
 wire \as2650.indirect_target[10] ;
 wire \as2650.indirect_target[11] ;
 wire \as2650.indirect_target[12] ;
 wire \as2650.indirect_target[13] ;
 wire \as2650.indirect_target[14] ;
 wire \as2650.indirect_target[15] ;
 wire \as2650.indirect_target[1] ;
 wire \as2650.indirect_target[2] ;
 wire \as2650.indirect_target[3] ;
 wire \as2650.indirect_target[4] ;
 wire \as2650.indirect_target[5] ;
 wire \as2650.indirect_target[6] ;
 wire \as2650.indirect_target[7] ;
 wire \as2650.indirect_target[8] ;
 wire \as2650.indirect_target[9] ;
 wire \as2650.insin[0] ;
 wire \as2650.insin[1] ;
 wire \as2650.insin[2] ;
 wire \as2650.insin[3] ;
 wire \as2650.insin[4] ;
 wire \as2650.insin[5] ;
 wire \as2650.insin[6] ;
 wire \as2650.insin[7] ;
 wire \as2650.instruction_args_latch[0] ;
 wire \as2650.instruction_args_latch[10] ;
 wire \as2650.instruction_args_latch[11] ;
 wire \as2650.instruction_args_latch[12] ;
 wire \as2650.instruction_args_latch[13] ;
 wire \as2650.instruction_args_latch[14] ;
 wire \as2650.instruction_args_latch[15] ;
 wire \as2650.instruction_args_latch[1] ;
 wire \as2650.instruction_args_latch[2] ;
 wire \as2650.instruction_args_latch[3] ;
 wire \as2650.instruction_args_latch[4] ;
 wire \as2650.instruction_args_latch[5] ;
 wire \as2650.instruction_args_latch[6] ;
 wire \as2650.instruction_args_latch[7] ;
 wire \as2650.instruction_args_latch[8] ;
 wire \as2650.instruction_args_latch[9] ;
 wire \as2650.io_bus_we ;
 wire \as2650.irqs_latch[1] ;
 wire \as2650.irqs_latch[2] ;
 wire \as2650.irqs_latch[3] ;
 wire \as2650.irqs_latch[4] ;
 wire \as2650.irqs_latch[5] ;
 wire \as2650.irqs_latch[6] ;
 wire \as2650.irqs_latch[7] ;
 wire \as2650.is_interrupt_cycle ;
 wire \as2650.ivectors_base[0] ;
 wire \as2650.ivectors_base[10] ;
 wire \as2650.ivectors_base[11] ;
 wire \as2650.ivectors_base[1] ;
 wire \as2650.ivectors_base[2] ;
 wire \as2650.ivectors_base[3] ;
 wire \as2650.ivectors_base[4] ;
 wire \as2650.ivectors_base[5] ;
 wire \as2650.ivectors_base[6] ;
 wire \as2650.ivectors_base[7] ;
 wire \as2650.ivectors_base[8] ;
 wire \as2650.ivectors_base[9] ;
 wire \as2650.page_reg[0] ;
 wire \as2650.page_reg[1] ;
 wire \as2650.page_reg[2] ;
 wire \as2650.regs[0][0] ;
 wire \as2650.regs[0][1] ;
 wire \as2650.regs[0][2] ;
 wire \as2650.regs[0][3] ;
 wire \as2650.regs[0][4] ;
 wire \as2650.regs[0][5] ;
 wire \as2650.regs[0][6] ;
 wire \as2650.regs[0][7] ;
 wire \as2650.regs[1][0] ;
 wire \as2650.regs[1][1] ;
 wire \as2650.regs[1][2] ;
 wire \as2650.regs[1][3] ;
 wire \as2650.regs[1][4] ;
 wire \as2650.regs[1][5] ;
 wire \as2650.regs[1][6] ;
 wire \as2650.regs[1][7] ;
 wire \as2650.regs[2][0] ;
 wire \as2650.regs[2][1] ;
 wire \as2650.regs[2][2] ;
 wire \as2650.regs[2][3] ;
 wire \as2650.regs[2][4] ;
 wire \as2650.regs[2][5] ;
 wire \as2650.regs[2][6] ;
 wire \as2650.regs[2][7] ;
 wire \as2650.regs[3][0] ;
 wire \as2650.regs[3][1] ;
 wire \as2650.regs[3][2] ;
 wire \as2650.regs[3][3] ;
 wire \as2650.regs[3][4] ;
 wire \as2650.regs[3][5] ;
 wire \as2650.regs[3][6] ;
 wire \as2650.regs[3][7] ;
 wire \as2650.regs[4][0] ;
 wire \as2650.regs[4][1] ;
 wire \as2650.regs[4][2] ;
 wire \as2650.regs[4][3] ;
 wire \as2650.regs[4][4] ;
 wire \as2650.regs[4][5] ;
 wire \as2650.regs[4][6] ;
 wire \as2650.regs[4][7] ;
 wire \as2650.regs[5][0] ;
 wire \as2650.regs[5][1] ;
 wire \as2650.regs[5][2] ;
 wire \as2650.regs[5][3] ;
 wire \as2650.regs[5][4] ;
 wire \as2650.regs[5][5] ;
 wire \as2650.regs[5][6] ;
 wire \as2650.regs[5][7] ;
 wire \as2650.regs[6][0] ;
 wire \as2650.regs[6][1] ;
 wire \as2650.regs[6][2] ;
 wire \as2650.regs[6][3] ;
 wire \as2650.regs[6][4] ;
 wire \as2650.regs[6][5] ;
 wire \as2650.regs[6][6] ;
 wire \as2650.regs[6][7] ;
 wire \as2650.regs[7][0] ;
 wire \as2650.regs[7][1] ;
 wire \as2650.regs[7][2] ;
 wire \as2650.regs[7][3] ;
 wire \as2650.regs[7][4] ;
 wire \as2650.regs[7][5] ;
 wire \as2650.regs[7][6] ;
 wire \as2650.regs[7][7] ;
 wire \as2650.relative_cyc ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][15] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[10][0] ;
 wire \as2650.stack[10][10] ;
 wire \as2650.stack[10][11] ;
 wire \as2650.stack[10][12] ;
 wire \as2650.stack[10][13] ;
 wire \as2650.stack[10][14] ;
 wire \as2650.stack[10][15] ;
 wire \as2650.stack[10][1] ;
 wire \as2650.stack[10][2] ;
 wire \as2650.stack[10][3] ;
 wire \as2650.stack[10][4] ;
 wire \as2650.stack[10][5] ;
 wire \as2650.stack[10][6] ;
 wire \as2650.stack[10][7] ;
 wire \as2650.stack[10][8] ;
 wire \as2650.stack[10][9] ;
 wire \as2650.stack[11][0] ;
 wire \as2650.stack[11][10] ;
 wire \as2650.stack[11][11] ;
 wire \as2650.stack[11][12] ;
 wire \as2650.stack[11][13] ;
 wire \as2650.stack[11][14] ;
 wire \as2650.stack[11][15] ;
 wire \as2650.stack[11][1] ;
 wire \as2650.stack[11][2] ;
 wire \as2650.stack[11][3] ;
 wire \as2650.stack[11][4] ;
 wire \as2650.stack[11][5] ;
 wire \as2650.stack[11][6] ;
 wire \as2650.stack[11][7] ;
 wire \as2650.stack[11][8] ;
 wire \as2650.stack[11][9] ;
 wire \as2650.stack[12][0] ;
 wire \as2650.stack[12][10] ;
 wire \as2650.stack[12][11] ;
 wire \as2650.stack[12][12] ;
 wire \as2650.stack[12][13] ;
 wire \as2650.stack[12][14] ;
 wire \as2650.stack[12][15] ;
 wire \as2650.stack[12][1] ;
 wire \as2650.stack[12][2] ;
 wire \as2650.stack[12][3] ;
 wire \as2650.stack[12][4] ;
 wire \as2650.stack[12][5] ;
 wire \as2650.stack[12][6] ;
 wire \as2650.stack[12][7] ;
 wire \as2650.stack[12][8] ;
 wire \as2650.stack[12][9] ;
 wire \as2650.stack[13][0] ;
 wire \as2650.stack[13][10] ;
 wire \as2650.stack[13][11] ;
 wire \as2650.stack[13][12] ;
 wire \as2650.stack[13][13] ;
 wire \as2650.stack[13][14] ;
 wire \as2650.stack[13][15] ;
 wire \as2650.stack[13][1] ;
 wire \as2650.stack[13][2] ;
 wire \as2650.stack[13][3] ;
 wire \as2650.stack[13][4] ;
 wire \as2650.stack[13][5] ;
 wire \as2650.stack[13][6] ;
 wire \as2650.stack[13][7] ;
 wire \as2650.stack[13][8] ;
 wire \as2650.stack[13][9] ;
 wire \as2650.stack[14][0] ;
 wire \as2650.stack[14][10] ;
 wire \as2650.stack[14][11] ;
 wire \as2650.stack[14][12] ;
 wire \as2650.stack[14][13] ;
 wire \as2650.stack[14][14] ;
 wire \as2650.stack[14][15] ;
 wire \as2650.stack[14][1] ;
 wire \as2650.stack[14][2] ;
 wire \as2650.stack[14][3] ;
 wire \as2650.stack[14][4] ;
 wire \as2650.stack[14][5] ;
 wire \as2650.stack[14][6] ;
 wire \as2650.stack[14][7] ;
 wire \as2650.stack[14][8] ;
 wire \as2650.stack[14][9] ;
 wire \as2650.stack[15][0] ;
 wire \as2650.stack[15][10] ;
 wire \as2650.stack[15][11] ;
 wire \as2650.stack[15][12] ;
 wire \as2650.stack[15][13] ;
 wire \as2650.stack[15][14] ;
 wire \as2650.stack[15][15] ;
 wire \as2650.stack[15][1] ;
 wire \as2650.stack[15][2] ;
 wire \as2650.stack[15][3] ;
 wire \as2650.stack[15][4] ;
 wire \as2650.stack[15][5] ;
 wire \as2650.stack[15][6] ;
 wire \as2650.stack[15][7] ;
 wire \as2650.stack[15][8] ;
 wire \as2650.stack[15][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][15] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][15] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][15] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][15] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][15] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][15] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][15] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack[8][0] ;
 wire \as2650.stack[8][10] ;
 wire \as2650.stack[8][11] ;
 wire \as2650.stack[8][12] ;
 wire \as2650.stack[8][13] ;
 wire \as2650.stack[8][14] ;
 wire \as2650.stack[8][15] ;
 wire \as2650.stack[8][1] ;
 wire \as2650.stack[8][2] ;
 wire \as2650.stack[8][3] ;
 wire \as2650.stack[8][4] ;
 wire \as2650.stack[8][5] ;
 wire \as2650.stack[8][6] ;
 wire \as2650.stack[8][7] ;
 wire \as2650.stack[8][8] ;
 wire \as2650.stack[8][9] ;
 wire \as2650.stack[9][0] ;
 wire \as2650.stack[9][10] ;
 wire \as2650.stack[9][11] ;
 wire \as2650.stack[9][12] ;
 wire \as2650.stack[9][13] ;
 wire \as2650.stack[9][14] ;
 wire \as2650.stack[9][15] ;
 wire \as2650.stack[9][1] ;
 wire \as2650.stack[9][2] ;
 wire \as2650.stack[9][3] ;
 wire \as2650.stack[9][4] ;
 wire \as2650.stack[9][5] ;
 wire \as2650.stack[9][6] ;
 wire \as2650.stack[9][7] ;
 wire \as2650.stack[9][8] ;
 wire \as2650.stack[9][9] ;
 wire \as2650.trap ;
 wire \as2650.warmup[0] ;
 wire \as2650.warmup[1] ;
 wire \as2650.wb_hidden_rom_enable ;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \wb_counter[0] ;
 wire \wb_counter[10] ;
 wire \wb_counter[11] ;
 wire \wb_counter[12] ;
 wire \wb_counter[13] ;
 wire \wb_counter[14] ;
 wire \wb_counter[15] ;
 wire \wb_counter[16] ;
 wire \wb_counter[17] ;
 wire \wb_counter[18] ;
 wire \wb_counter[19] ;
 wire \wb_counter[1] ;
 wire \wb_counter[20] ;
 wire \wb_counter[21] ;
 wire \wb_counter[22] ;
 wire \wb_counter[23] ;
 wire \wb_counter[24] ;
 wire \wb_counter[25] ;
 wire \wb_counter[26] ;
 wire \wb_counter[27] ;
 wire \wb_counter[28] ;
 wire \wb_counter[29] ;
 wire \wb_counter[2] ;
 wire \wb_counter[30] ;
 wire \wb_counter[31] ;
 wire \wb_counter[3] ;
 wire \wb_counter[4] ;
 wire \wb_counter[5] ;
 wire \wb_counter[6] ;
 wire \wb_counter[7] ;
 wire \wb_counter[8] ;
 wire \wb_counter[9] ;
 wire wb_debug_carry;
 wire wb_debug_cc;
 wire wb_feedback_delay;
 wire wb_io3_test;
 wire wb_reset_override;
 wire wb_reset_override_en;
 wire \web_behavior[0] ;
 wire \web_behavior[1] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__A1 (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__A2 (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__A1 (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05665__I (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05667__I (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05670__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__I (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__A2 (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05675__I (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05678__A3 (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05678__A4 (.I(\as2650.is_interrupt_cycle ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05680__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__A1 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05683__I (.I(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05686__A2 (.I(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05686__B1 (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05687__A2 (.I(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05687__B1 (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05688__I (.I(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05691__B2 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05692__B2 (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05694__A1 (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05694__A2 (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05695__A1 (.I(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05696__A2 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05697__B1 (.I(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05697__B2 (.I(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__A2 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__B1 (.I(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__B2 (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05701__A1 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05701__A2 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05703__A2 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05703__B2 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05704__B2 (.I(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05707__A1 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05707__A3 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__A2 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__B1 (.I(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05709__A3 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05711__A1 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05711__A2 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05711__A3 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__A1 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05713__A1 (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05713__A2 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05716__B2 (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05717__A1 (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05717__A2 (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05717__A4 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05719__A1 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05721__B2 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05731__A2 (.I(\as2650.cpu_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__A1 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__A2 (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__A1 (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__A2 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__A3 (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__A1 (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__A2 (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__A3 (.I(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05737__I1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05737__S (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__A2 (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05741__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05741__A2 (.I(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__I (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__A1 (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__A2 (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__A3 (.I(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__B (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__A1 (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__A3 (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__A4 (.I(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05749__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05751__A2 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05751__A3 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__I (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05755__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__I (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__I (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__I (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__I (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A1 (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__I (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05766__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__S (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__I (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__I (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__A2 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__A2 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__I (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__A1 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__A1 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__I (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__I0 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__I1 (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__I (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__A1 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__A2 (.I(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__B2 (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__C (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__I (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__A1 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__A1 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__I (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05800__S (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__I0 (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__I1 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__A1 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__I (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05808__I (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__A1 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__I0 (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__I1 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__S (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__A4 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__A1 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__A1 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__I0 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__I1 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__A1 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__A1 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A1 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__I0 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__S (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__I (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A1 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__A1 (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05836__A2 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__A1 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__A2 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__A2 (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__A1 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__A1 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__S (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__I0 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__I1 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__A1 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__A1 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__I (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05853__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05854__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__A2 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A2 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A1 (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A2 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__A2 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__B (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A2 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A3 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__S (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__I (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__S (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__I0 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__I1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__A1 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__I0 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A2 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__A2 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__A1 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__A1 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__S (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__I (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__A2 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__A2 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__I (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__I0 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__I1 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__I (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__A1 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__A2 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__A2 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__B (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A2 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A3 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__I (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A1 (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__A2 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__A2 (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A1 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__I (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__S (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__I (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A2 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__I0 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__I1 (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A2 (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A2 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__C (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__A2 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A1 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A2 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__B (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A1 (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__A2 (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__A2 (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A1 (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__I (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__S (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__I (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A2 (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__A2 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__I0 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__I1 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__A2 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__A1 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__A2 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A1 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A2 (.I(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A4 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A2 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A3 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__B (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__A2 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__B (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05984__A2 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__A2 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__A1 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__A1 (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__A2 (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__I (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__A1 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__A3 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__I (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__A1 (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A1 (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__A1 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__A2 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__I (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A1 (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A3 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A1 (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__A1 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A1 (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A2 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__A1 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__A1 (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__A2 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__A2 (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__A3 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__A4 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__I (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A1 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__A1 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__I (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A2 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__B1 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__B2 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__A2 (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__A1 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__A3 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A1 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A2 (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__A2 (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A2 (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__I (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A2 (.I(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__B1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__B2 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__A2 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__A2 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A2 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A2 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__A1 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A1 (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__A1 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__A3 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__A3 (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A1 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A1 (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A3 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__A1 (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__A3 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A2 (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A1 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A1 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A3 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A1 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A3 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__A1 (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__A1 (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__A3 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__A3 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__I (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__I (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__I (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A1 (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A2 (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A4 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__A2 (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__I (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__I (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__A2 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__A2 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A2 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A2 (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A2 (.I(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__I (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__I (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__I (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__I (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__I (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__I (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__I (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__I (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__I (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__I (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__I (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__I (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__I (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__I (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__I (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A2 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__A1 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__A2 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__A2 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__A2 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A1 (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__A2 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__A2 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__A4 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A2 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A1 (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A2 (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__A2 (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__A2 (.I(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__B1 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__B2 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A1 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__B (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A2 (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__B2 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__C (.I(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A1 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A2 (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__A1 (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__A2 (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__A2 (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__A2 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A2 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A1 (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A2 (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__A1 (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__A2 (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A1 (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A2 (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__A1 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__I (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__I (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A1 (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__A2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__A3 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A3 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A4 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A2 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__B (.I(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__I (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A3 (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06189__I (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__I (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A2 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A2 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__I1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__I0 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__I1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__I1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__S (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__I1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__A2 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__A2 (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A2 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__I (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__A1 (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__A3 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A1 (.I(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A2 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__A2 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__I (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A1 (.I(\as2650.insin[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A1 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A2 (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A2 (.I(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__A1 (.I(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A1 (.I(\as2650.insin[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A2 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A1 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A2 (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__A2 (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A2 (.I(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A2 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A2 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A3 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A1 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__I (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A1 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A2 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__B (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A2 (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__I (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__I (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A2 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A1 (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A2 (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__I (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A2 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__I (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A3 (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__I (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__I (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A1 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A2 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__I (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__I (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A2 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__A1 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A1 (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A2 (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A1 (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__I (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A2 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A3 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__I (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__I (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__I (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A1 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A1 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__B (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A2 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__I (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__I (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__I (.I(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__I (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__I (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A2 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__A1 (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__A2 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__A2 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__I (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A1 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A2 (.I(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A1 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A3 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__I (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__I (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__I (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__A2 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__I (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A1 (.I(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A2 (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A4 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__A2 (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__I (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__B (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__B1 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A2 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A2 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__A2 (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A2 (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__I (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__I (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A1 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A2 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A1 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__A1 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__B (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A2 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A1 (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A2 (.I(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A2 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A3 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__A2 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__A3 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A1 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A2 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A1 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A2 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A1 (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A1 (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__I (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__I (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A1 (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__I (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__I (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__I (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__I0 (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__I1 (.I(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__S (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__I (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__I0 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A1 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A2 (.I(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__A1 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__A2 (.I(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__I (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A2 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__I (.I(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__I (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A1 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A3 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A4 (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__A1 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__A1 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A1 (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A2 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__B2 (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__A1 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__I (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__I (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A1 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A2 (.I(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A1 (.I(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__B1 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__I (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__I (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A1 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A1 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A1 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__B1 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__I (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__A1 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__I (.I(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A1 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__A1 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__B1 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__I0 (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__S (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__S (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__I (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__I (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__A1 (.I(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__A2 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__A1 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__B1 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A1 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__B (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__I (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06480__A1 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06480__A2 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A2 (.I(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A3 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A2 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A3 (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__B1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A1 (.I(\as2650.debug_psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A2 (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A1 (.I(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A2 (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__B (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__C (.I(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__A1 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__A1 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A2 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A3 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A2 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A3 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__I (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__I (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__I (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__A2 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A2 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__I (.I(\as2650.is_interrupt_cycle ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__I (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A2 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A1 (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__I (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__A1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__A1 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__A3 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__I (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__I (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__I (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__A1 (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__A2 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__A3 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__A1 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__A2 (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__I (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__A1 (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__A2 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__B (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__I (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__A1 (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__A2 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__A1 (.I(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A1 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A2 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A3 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__I (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__C (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__B2 (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__A2 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__A2 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__A3 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A2 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A2 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A3 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A3 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A2 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__A1 (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__I (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__I (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A1 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A4 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__I (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__I (.I(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__B (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__I (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__C (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__I (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__I (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__I (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__I (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__I (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__I (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__I (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A1 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A2 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__B (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A1 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__C (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__I (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__I (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__I (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__A2 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A2 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A3 (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A4 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A1 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A3 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__I (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A2 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__B2 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__I (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A2 (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__I (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A2 (.I(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A2 (.I(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__B (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__I (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__I (.I(\as2650.debug_psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__I (.I(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A3 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A2 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A2 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__I (.I(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__A1 (.I(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__A3 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__A2 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__I (.I(\as2650.debug_psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__I (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__I (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__A2 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__I (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__I (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__I (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__I (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__I (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A1 (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A2 (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A2 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__A4 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__I (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A1 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__A1 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A2 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__A1 (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__I (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__I (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__I (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__I (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A2 (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__A2 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A1 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A1 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__B (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__A1 (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__I (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__I (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__I0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__I1 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__S (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A1 (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A2 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A2 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__A1 (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__I (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__I (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__I0 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__I (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A1 (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A2 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__B (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A1 (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__I (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__I0 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__I1 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__S (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__I (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A2 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__B (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__A1 (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A1 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__I (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A2 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A2 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__I (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A1 (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__B (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A1 (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__I (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__A2 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A1 (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A2 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__B (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A1 (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__I (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__I (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A1 (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A2 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A2 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__I (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__A1 (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__B (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A1 (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A1 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__I (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A2 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A2 (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__I (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A1 (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__B (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A1 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__I (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__I (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A2 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__I (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__I (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A2 (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A3 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__I (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__I (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__I (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__A1 (.I(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__I (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A1 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A2 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__I (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__I (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__B (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A1 (.I(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A2 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A1 (.I(net427));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A2 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A3 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__I (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__I0 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__I1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__I0 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__I1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__I0 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__I1 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__I0 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__I1 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__I (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__I0 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__I1 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__I0 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__I1 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__I0 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__I1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__I0 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__I1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__I (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__I0 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__I1 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__I0 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__I1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__I0 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__I1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__I0 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__I1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__I (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__I0 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__I1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__I0 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__I1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__I0 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__I1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__I0 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__I1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__I (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__I1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__I0 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__I1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__I1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__I1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__I (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__I1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__I0 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__I1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__I0 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__I1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__I0 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__I1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__I (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__I0 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__I1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__I0 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__I1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__I0 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__I1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__I0 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__I1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__I (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__I0 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__I1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__S (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__I0 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__I1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__S (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__I0 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__I1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__S (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__I0 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__I1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__S (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__I (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__I (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A1 (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__C (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A2 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A3 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A4 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A2 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I0 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__S (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I0 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__S (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__I0 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__I1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__S (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__I (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A2 (.I(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A1 (.I(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A2 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__I (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__I (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A2 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__B1 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__B2 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A2 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A1 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A1 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__C (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__A1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__A2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__I (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__I (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__B (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__C (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A2 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A1 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__A1 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__C (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A1 (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A2 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__B (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__C (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A2 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A1 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__C (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__I (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__I (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A1 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A2 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__I (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__I (.I(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__I (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A1 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__B2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__C (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A1 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A2 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A1 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A1 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__I (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__I (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__B (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__B2 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__C (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A1 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A1 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A1 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A2 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__B (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__I (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__B (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__I (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A1 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A2 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__B (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A1 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__I (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__I (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__I (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__I (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__I (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__I (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07056__A2 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__I (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A2 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A2 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__I (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A2 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__I (.I(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A2 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__I (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A2 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__B (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__I (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A2 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A2 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__B (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A1 (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A2 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__B (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__I (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A3 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__I (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__A1 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__I (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__C (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__A1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__I (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__C (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__I (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__B (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__C (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__I (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__C (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__I (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__I (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__C (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__I (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__C (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__C (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__B (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__I (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__B1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__I (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__I (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__I (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A1 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__B (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A1 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__I (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__B (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A1 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__I (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__C (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__I (.I(net287));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A2 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__B (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A1 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__B (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A2 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__C (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A2 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__B (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__B (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A2 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__C (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A2 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A2 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__C (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__B (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A2 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__C (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A2 (.I(net441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A2 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A4 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__I (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__I (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__I (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__B (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A1 (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__C (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__B (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A2 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__A2 (.I(net437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__C (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__I (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__I (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__I (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A2 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A1 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A1 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__I (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__A2 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__C (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__I (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A1 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__I (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__I (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__I (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__I (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__I (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A1 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A1 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A1 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__I (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A1 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__I (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__I (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07332__I (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__I (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__I (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__I (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__I (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__I (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__I (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__I (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__B (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__B (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__B (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__B (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A1 (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A1 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__B (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A1 (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A2 (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A1 (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A2 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A1 (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__B (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__I (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A1 (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A2 (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__A1 (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__A2 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A1 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A1 (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__B (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A1 (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A1 (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A2 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A1 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A1 (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__B (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__I (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A1 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A2 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__B (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__I (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__I (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A1 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A2 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A2 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A3 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A2 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A2 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__I (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A1 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A2 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A3 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A2 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__I (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A2 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__B (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__I (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A2 (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__I (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__I (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__I (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__I (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A1 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A2 (.I(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__I (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__I (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__I (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__I (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__I (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__I (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__I (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__I (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__I (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__I (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__I (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__B2 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__A1 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__I (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__I (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__I (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__C (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A1 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__I (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__I (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__I (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A1 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__I (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__C (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A1 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__I (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__I (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__I (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__S (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__I (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__I (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A1 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__B2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__I (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__I (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__I (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A1 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A2 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A3 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__A2 (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__I (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__I (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__I (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__I (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A2 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A3 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__I (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A1 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A2 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__I (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A2 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__B (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__C (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__I (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__I (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__I (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__I (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__I (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__B1 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__B2 (.I(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__C (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__I (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__I (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__I (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__I (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__B1 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__B2 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__C (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__I (.I(\as2650.is_interrupt_cycle ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__I (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__I (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__I (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__I (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__I (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A1 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A2 (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__I0 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__I1 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__I (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__I (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A2 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__B2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__B (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__I (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__I (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__I (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__I (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__I (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A2 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__B2 (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__B (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__I (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__I (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__I (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__I (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A2 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__B1 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__B2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__C (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__I (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__I (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__I (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__I (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(\as2650.insin[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__B1 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__B2 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__C (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A2 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__I (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A1 (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__I (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__A2 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A1 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A4 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__I (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A2 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__A2 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__I (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__B2 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__A2 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__A2 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__B (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A2 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A1 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A2 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A3 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__I (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A1 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A3 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__B (.I(\as2650.cpu_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__C (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A2 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__I (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__B (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__I (.I(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__I (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__I (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__I (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A2 (.I(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A1 (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A3 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__I (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__B2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A1 (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__B2 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__I (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__B2 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A1 (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__I (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__I (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A2 (.I(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__A1 (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A1 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A1 (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A1 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__B2 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__A1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__B1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__B2 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__I (.I(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__A3 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A1 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__B2 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__B1 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__B2 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__B2 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__A2 (.I(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__I (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__I (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__I (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__I (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A1 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A1 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A2 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__B1 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__B2 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__B1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__B2 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__C (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A1 (.I(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A2 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__I (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__I (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__I (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__I (.I(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A1 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__I (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A1 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A1 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A1 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__B2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A1 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__B1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__B2 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__I (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A1 (.I(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A2 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__I (.I(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__I (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__I (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A2 (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A2 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A3 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A1 (.I(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A1 (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A1 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A1 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__A1 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A2 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__B2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__B1 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__B2 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__I (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A1 (.I(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__I (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__I (.I(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A2 (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__B (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__I (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A1 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__A2 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A2 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__B2 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__B1 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__B2 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A1 (.I(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__I (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A2 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__B1 (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__B2 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A1 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__B1 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__B2 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A1 (.I(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__I (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A1 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A2 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__I (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A1 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__I (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A1 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__B1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__B2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__C (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__A1 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__A2 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A1 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__B (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A2 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__I (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A1 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__C (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__I (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__I (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__C (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__I (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__I (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A2 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A1 (.I(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__I (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A1 (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__I (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A2 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A3 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__I (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__I (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__I (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__C (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__C (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A2 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A3 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A1 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__C (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__C (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__I (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__B2 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__C (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__I (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__I (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A1 (.I(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__B (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A2 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__I (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__I (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__B (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__C (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A2 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A4 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A1 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A3 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__I (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A2 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__B (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__C (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__A1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A1 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A3 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__B (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__C (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A2 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A3 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A2 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__B1 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A1 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__B (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__I (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__I (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A1 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A1 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A3 (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__A2 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__B (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__I (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A1 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A2 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__B (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__I (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__B (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A1 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A1 (.I(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__I (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__I (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A2 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A3 (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A1 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__I (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__I (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A2 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A3 (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A1 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A2 (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A3 (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A1 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__I (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__I (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__I (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A2 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__I (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A2 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__B1 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__I (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A2 (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A2 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A1 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__B2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__I (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A1 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A2 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__B1 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__I (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A2 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__I (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__I (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A2 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__B1 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__B1 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A1 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__I (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__I (.I(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__I (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__I (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A1 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A2 (.I(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__B1 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A2 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A3 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__B1 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__I (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A2 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A3 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__I (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__I (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A1 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A2 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__B1 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A2 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A3 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A3 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A2 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__B2 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__B2 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__I (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A2 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A2 (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__B2 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__B2 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__I (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__B2 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A2 (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__B2 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A3 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__B2 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A3 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A3 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__B2 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A1 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__B1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A3 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A1 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A2 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A1 (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A2 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__I (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__I (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__I (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A1 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A2 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A1 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A2 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A1 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A1 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A2 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__A1 (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A1 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A2 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A3 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A4 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A2 (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__I (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A1 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A2 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A1 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A1 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A2 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A1 (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A2 (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__A1 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A1 (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__B (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A2 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A3 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A1 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A2 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A3 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__I (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__I (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A2 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A3 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A1 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A1 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__C (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__I (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__I (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__I (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__I (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__I (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__I (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__I (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A1 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A1 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__I (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__I (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__I (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__I (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__I (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__I (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__I (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__C (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__I (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__I (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__I (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__I (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__I (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__I (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A2 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__C (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A1 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__C (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__I (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__I (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__A1 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A2 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__C (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__I (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__S (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A1 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A1 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__B (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__B (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__I (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A1 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__C (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A1 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__C (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A1 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A2 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__C (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__I (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__C (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__I (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__I (.I(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A1 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__C (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__S (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__I (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__B (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__I (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A2 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A3 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A4 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A1 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__I (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A1 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A4 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A1 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A1 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A1 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A1 (.I(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A2 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__B (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A1 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A1 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A1 (.I(\as2650.insin[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A2 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__B (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A3 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__I (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__A1 (.I(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__B (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__I (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A1 (.I(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__B (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A1 (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__I (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__I (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A1 (.I(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__I (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A1 (.I(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__I (.I(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__I (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__A1 (.I(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A1 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__I (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__A1 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A1 (.I(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__I (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A1 (.I(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A1 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__I (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__I (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__I (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__B (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__B (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A1 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A1 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A2 (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A1 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__B1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__C (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__B1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__B1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__C (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A2 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__B1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__S (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A3 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__B (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__I (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A3 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__B (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A2 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A3 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__I (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A1 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__B (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A1 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A2 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A1 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__I (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__C (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__I (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A2 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A2 (.I(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A2 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A1 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__I (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__B2 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__C (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__I (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__I (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A1 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__C (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__I (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A1 (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__B (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__I (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A2 (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__C (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__I (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__I (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A2 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__B2 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__C (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A2 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A2 (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__C (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A2 (.I(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A2 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A2 (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__B2 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__C (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__S (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__I (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A2 (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A3 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__B1 (.I(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A2 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A1 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__B2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A1 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__C (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__A1 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__B (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__C (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__I (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A1 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__B (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__I (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__C (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A2 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__C (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__S (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__A1 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__B1 (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__B (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A1 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A2 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__B (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A2 (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__B1 (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__B2 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A1 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__B (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__I (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A2 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__B1 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__C (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A2 (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A2 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__B (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A2 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__B1 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__B2 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__C (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__B (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__B2 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__C (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A1 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A2 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__B (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A2 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__B1 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__B2 (.I(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__S (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A1 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__B1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__B2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A2 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__I (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__I (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__B2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__I (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__I (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__B1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__B2 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__C (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A1 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__I (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__I (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A1 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__B (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__B1 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__C (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__B (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A2 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A2 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__B (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A2 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__B1 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__C (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A2 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__B (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A2 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__B2 (.I(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__S (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__B1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__B (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A2 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__I (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__C (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A1 (.I(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__C (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__I (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A3 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A1 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__B (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__B1 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__B2 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__C (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__B (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__C (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A1 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__B (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__B1 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__C (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A1 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A1 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A2 (.I(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__B (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A1 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__B1 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__B2 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__C (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__S (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__B1 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__B (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__I (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__A1 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__C (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A1 (.I(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A1 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A2 (.I(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__C (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__I (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A1 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__I (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A2 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__B2 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__C (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__C (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__S (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__B1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__B (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A1 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__B2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__A1 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__B2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__A1 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A1 (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A2 (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__B2 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__C (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A2 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__I (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A1 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__I (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__B1 (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__C (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A2 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__B1 (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__C (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A2 (.I(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__B2 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__C (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__S (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__B1 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__B2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__B (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__B2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__C (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A1 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__C (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__A2 (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A1 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__B (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__I (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__B1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__B (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__I (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__C (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__B (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__B1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__C (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__B (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__C (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__B1 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__S (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__B1 (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__B2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__C (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A1 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A2 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__B2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A1 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__A1 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A2 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A1 (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__B2 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__C (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__I (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A1 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__A1 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__B (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__B (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__I (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__I (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__I (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__B1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__C (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__B (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__B (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__B1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__C (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__S (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__B1 (.I(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A1 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A1 (.I(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A1 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A2 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A2 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A1 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A2 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__B2 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__C (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A1 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A2 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__B (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A1 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__B2 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A1 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A2 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__A1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__B (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__B1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__C (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A1 (.I(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__B (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A2 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__B1 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__C (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A2 (.I(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__B (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__B1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A1 (.I(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A1 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__B (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__B1 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__C (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__S (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__B1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__B2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__C (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A1 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A1 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A3 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A4 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__I (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__I (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A1 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__B (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__I (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__B1 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__C (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__B (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__B1 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__C (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A1 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__B1 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__C (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__B (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__B1 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__C (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__I1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__S (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__B1 (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A1 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A1 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A2 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__C (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A2 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A1 (.I(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__B2 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__B (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__I (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A2 (.I(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__I (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__B2 (.I(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A1 (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__C (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__A1 (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__C (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__S (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__A1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__B1 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A2 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A1 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__B2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A1 (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A1 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A1 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__B2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A2 (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A1 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__I (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A2 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__I (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A1 (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A2 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A2 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__B (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__C (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__I (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__I (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A2 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A2 (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A1 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A2 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__I (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A1 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A2 (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A2 (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A2 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A1 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A2 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A1 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__I0 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__I1 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A2 (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__I (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A2 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__I0 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__I1 (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A2 (.I(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A1 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A2 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A2 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A2 (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__B (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A2 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__I (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__C (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__I (.I(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A2 (.I(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A2 (.I(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__I (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A2 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A2 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A3 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A3 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__B2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__I (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A1 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A3 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A2 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__B (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A1 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A2 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__B (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A2 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__I (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__I (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__I (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A2 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__I (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A2 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__B2 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__I (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A3 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A2 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A3 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A2 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A2 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__B (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__I (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A2 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__I (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A2 (.I(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__B1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__B2 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__B2 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A1 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A2 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__I (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A2 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A3 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__I (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__B (.I(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A2 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A2 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A3 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__I (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A1 (.I(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A2 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__B1 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__C (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__I (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A2 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A1 (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A2 (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A1 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__C (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A2 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__B (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A1 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__B (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A1 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A2 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A3 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A2 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__I (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__B (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A2 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A2 (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__B1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__B2 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__B2 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A1 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A2 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__B (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__I (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__B (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__B (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A1 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__C2 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A1 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A1 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__B1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A1 (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__I (.I(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__B2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A1 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A2 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A2 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__C (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__S1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A2 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__I2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__I3 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__I1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__S1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__I1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A3 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__I2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__I0 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__I2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__I3 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__I2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__I0 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A2 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A3 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A4 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A2 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__A2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A2 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__B1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__B2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A1 (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A2 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A2 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A2 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__B1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__B2 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A2 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__B1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__B2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A1 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__B1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__B2 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A1 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A2 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A3 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A2 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A1 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A1 (.I(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A2 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A3 (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A4 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A3 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A1 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A2 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A3 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A4 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__I (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A2 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__A1 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A1 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A1 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__I (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A1 (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A1 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__B2 (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__I (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A2 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A1 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A1 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A2 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__B1 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__B2 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A1 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A2 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A2 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A1 (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__B2 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A2 (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A1 (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__I (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A1 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A1 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A2 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A2 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A1 (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A2 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A1 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A2 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A2 (.I(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A2 (.I(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A1 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__B2 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__B2 (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A3 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A2 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__B2 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A2 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A3 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A4 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__I (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A2 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A2 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A4 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__B1 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A2 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A1 (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A2 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A1 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A1 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A2 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__A2 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__I (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A1 (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A1 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A2 (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__B (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__C (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A2 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__B1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__B2 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A3 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A1 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(\as2650.debug_psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__I (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__I (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A2 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A3 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A4 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A2 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A3 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A4 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__B (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A1 (.I(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A2 (.I(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__B1 (.I(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__C (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__B1 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__A1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__B2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__C (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__B1 (.I(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A2 (.I(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__C (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A2 (.I(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__C (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__B1 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A2 (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A3 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A4 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__C (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A2 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A1 (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A2 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__B1 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__B2 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__A2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__B1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__B2 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A2 (.I(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__B1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__B2 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A1 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A1 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A2 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A2 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__B2 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A1 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A2 (.I(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__B1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__B2 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A2 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A1 (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A3 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A1 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A2 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A3 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A2 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__B (.I(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A1 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__B2 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__B2 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A2 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A2 (.I(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__I (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__B1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__B2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__C1 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__C2 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__I (.I(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__B1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__B2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A2 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__B1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__B2 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A1 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__B (.I(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__B (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A1 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__I0 (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__I1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A2 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__B1 (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__B2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A1 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A2 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__B1 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__B2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A2 (.I(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09642__A1 (.I(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A1 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A1 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A2 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A1 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A1 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__B1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__B2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__B (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A3 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A2 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A3 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A2 (.I(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A3 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A4 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__B (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__B1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__B (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A2 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__B2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A2 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__B1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__B2 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A2 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__B1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__B2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A1 (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A1 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A2 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__B (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__C (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__I (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A1 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__I (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A2 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A2 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A1 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__B (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A2 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__C (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__I0 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A2 (.I(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A2 (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A2 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A2 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A2 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A3 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A1 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__B (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__I (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__B (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__I (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A1 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A2 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A1 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A2 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__B (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__B2 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A1 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A1 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__A1 (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__I (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A1 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A2 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A1 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A2 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A1 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A2 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A4 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A1 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A1 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A1 (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A2 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__I (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A2 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__A1 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A1 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A2 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__A3 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__B (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__B (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__C (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A2 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A1 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A1 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__A1 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A1 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A2 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__A1 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A3 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A1 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__A2 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A2 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__B (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A1 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A2 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A2 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A2 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A2 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A3 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__C (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A1 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__B2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__A1 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A1 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A3 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__B2 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__A1 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__B2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__B2 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__I1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__I1 (.I(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__I1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A2 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A1 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A2 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A2 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__B2 (.I(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A1 (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__I (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A2 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__B (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A2 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A2 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__B (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A2 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__I (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A2 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A2 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A2 (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A2 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__I (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A2 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__A2 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A2 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A2 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__I (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A2 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A2 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A2 (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A2 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A2 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A2 (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A1 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__I (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__I (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__B (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A1 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__B (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A1 (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A2 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A2 (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A2 (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__I (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A1 (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__B (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A2 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__B (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A1 (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__B (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A1 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A2 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A1 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__B (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A2 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__B (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__C (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A2 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__B (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A2 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__B (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__C (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A1 (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A2 (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__I (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A1 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A3 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A4 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A2 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A3 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A4 (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A2 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__B (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__I (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__I (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A3 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__A1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A2 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__I (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__I (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A2 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__A1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__A2 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__A1 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A1 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__I (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__I (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__I (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__I (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__I (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A1 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__B (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__I (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A2 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__I (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__I0 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A1 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__A2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__B (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__A1 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A2 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__B (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__I (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__I (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A1 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A2 (.I(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__B (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__I (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__I (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A2 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__I (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__I (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A3 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__I (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__I (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A1 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A1 (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__B (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__I (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A2 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A1 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__I0 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__B (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__I (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A2 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A1 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A1 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__B (.I(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__I (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A2 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A1 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__I (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__I0 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__I1 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__I (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__B (.I(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__I (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__I (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__I0 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__I1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A1 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__B (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__I (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__A1 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A1 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__A2 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__B (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__I (.I(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__I0 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__I1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__I (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__I (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__I0 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__I1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A1 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__A1 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__I (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__I (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A1 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__I (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A1 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__A1 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A1 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A2 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__B (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__I (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__I (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__I (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__I (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__I (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__I (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__I (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__I (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__A2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__B (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__I (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__I (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A1 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A1 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__I (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__I (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A2 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A2 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A2 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A2 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__I (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__I (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__I (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__I (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A2 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A2 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A2 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A2 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A2 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A2 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__A2 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A2 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__I (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__I (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A1 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__I (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__I (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A2 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A2 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A2 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__I (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__I (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__I (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__I (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A2 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A2 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__A2 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A2 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A2 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A2 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A2 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A2 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__I (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A1 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__I (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__I (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A2 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A2 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__I (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__A2 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__A2 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A2 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A2 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__I (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A2 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A2 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__I (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__I (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__I (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__I (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__I (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__I (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__I (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__I (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A1 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__I (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__I (.I(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__I (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__I (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__I (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__I (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A1 (.I(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__I (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A1 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A2 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A3 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__I (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__I (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A1 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__I (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A1 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__I (.I(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A1 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__I (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A2 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A1 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A1 (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__B (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A2 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__B2 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A3 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A1 (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__B (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A2 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A1 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A1 (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A2 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A4 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__I (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__I (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__I (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A1 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A1 (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A2 (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__I (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A2 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__I (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__B (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__I (.I(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__I (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__I (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A1 (.I(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A1 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A2 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__I (.I(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A2 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A3 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A2 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A3 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A2 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A3 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A3 (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__B (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A1 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A1 (.I(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A4 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A1 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A1 (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A2 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A4 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A2 (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A3 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A4 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__A2 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__B (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A1 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A1 (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A2 (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A4 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A2 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A2 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__A1 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A2 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A2 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A1 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A1 (.I(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A2 (.I(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__I (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__I (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__I (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__B2 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__B2 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A2 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A1 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A2 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A2 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__I (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A1 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A1 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__A2 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__I (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__I (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A1 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__B1 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A1 (.I(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A2 (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__I (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__I (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__I (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__I (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__A1 (.I(\as2650.debug_psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__A2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__I (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A2 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__B2 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A1 (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A1 (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__I (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A1 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A2 (.I(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__I (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__B1 (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A1 (.I(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A2 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__I (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__B (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__B1 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__B2 (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A1 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__B (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A1 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A2 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__I (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A1 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__C (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__I (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__A2 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A1 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__A1 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A1 (.I(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__A2 (.I(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__A1 (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__B1 (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__A1 (.I(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__A2 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__I (.I(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A1 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A2 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A1 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A2 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A1 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__C (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A1 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A1 (.I(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A2 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A2 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__A1 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__I0 (.I(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__I1 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__I (.I(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A1 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__B1 (.I(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A2 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__I (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A2 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__B1 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__B2 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A1 (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A1 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A1 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A1 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__C (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A1 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A1 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A2 (.I(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__I (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A1 (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__A1 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__B1 (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A1 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__A1 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__B1 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__B2 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__A1 (.I(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__A2 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__B (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A1 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A1 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A1 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A1 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__B (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A1 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__B (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A2 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__I0 (.I(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__I1 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__I (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__B1 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A2 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__I (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__B2 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__B1 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__B2 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__B (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10569__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__B (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__A1 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A2 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__B1 (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__C (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__A1 (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__A2 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A1 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A1 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A2 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__A1 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__I (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A1 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A1 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__B1 (.I(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__A1 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__I (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__I (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A2 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A2 (.I(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__A2 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A2 (.I(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A2 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A2 (.I(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__A2 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A2 (.I(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__I (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__I (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__I (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__I (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__A1 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__A1 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A1 (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__I (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__I (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A1 (.I(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A1 (.I(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A1 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A1 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__A1 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__I (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__I (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A2 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A2 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A2 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__A2 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__I (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__I (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A2 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__I (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__I (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A1 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__A1 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A1 (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__I (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__I (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A1 (.I(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__A1 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A2 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__I (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__I (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__I (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__I (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A1 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__I (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__I (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__A1 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A1 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__I (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__I (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A1 (.I(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A2 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A1 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A2 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A2 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__A2 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A1 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A1 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A1 (.I(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__A1 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A1 (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A1 (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__A1 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__A1 (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__A1 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__A1 (.I(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A1 (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__A1 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A1 (.I(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A3 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__I (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A2 (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__B1 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A1 (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__B1 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A1 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__B1 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A1 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__B1 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__I (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__I (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A2 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__I (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__I (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__I (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__I (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__I (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__I (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__I (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__I (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__I (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__I (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A1 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__I (.I(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A1 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__I (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A1 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__I (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__I (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__I (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A3 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__I (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A2 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A1 (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A1 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__A1 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__I (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A3 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__I (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A2 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A1 (.I(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A1 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__A1 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A1 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__I (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A1 (.I(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__A1 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A1 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__I (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A1 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A2 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__I (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__I (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__I (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__I (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A2 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A2 (.I(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__A2 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A2 (.I(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A2 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__A2 (.I(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__A2 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A2 (.I(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__I (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__I (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A1 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A1 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A1 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__I (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__I (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__I (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__I (.I(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__I (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__I (.I(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A2 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A2 (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A2 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A2 (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A2 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A2 (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A2 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A2 (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__I (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__I (.I(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A1 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A1 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__I (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__I (.I(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A2 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A2 (.I(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A2 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A2 (.I(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A2 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A2 (.I(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A2 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A2 (.I(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A1 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A3 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A4 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A2 (.I(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A2 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A2 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A2 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A2 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A1 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A2 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A2 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A1 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A1 (.I(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__B (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__I (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A1 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A2 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A1 (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__A2 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A2 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A2 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A1 (.I(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A1 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__B (.I(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A1 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__A1 (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__I (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A1 (.I(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A3 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__B2 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A2 (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A2 (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A2 (.I(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A1 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A1 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A1 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__A3 (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A1 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A2 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__A1 (.I(\as2650.chirpchar[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A1 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A1 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__I0 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A1 (.I(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A3 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__B2 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A2 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A1 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A1 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A1 (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A1 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A2 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__C (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__A1 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__A1 (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__A1 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__A2 (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__I (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__A1 (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__B2 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__A2 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__B (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__B1 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__C1 (.I(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__C2 (.I(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__A1 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__A2 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__I (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__I (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A1 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__I (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__I (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__I (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__I (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A1 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__A1 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__I (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__I (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A2 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A2 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__A2 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A2 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__A1 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__A2 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__I (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A3 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A1 (.I(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A2 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__A2 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A1 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A3 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A1 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__A1 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A1 (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__A1 (.I(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__A2 (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A3 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__A1 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__A2 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__A3 (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A1 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A1 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A1 (.I(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A3 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A1 (.I(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__A1 (.I(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__A3 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A1 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A1 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A1 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A1 (.I(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A3 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A1 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__A1 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A1 (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A2 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A3 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A2 (.I(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A1 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A3 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A3 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__I (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A2 (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A1 (.I(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__A1 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A1 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A1 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__I (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A1 (.I(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A1 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A1 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__I (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__I (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__I (.I(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__I (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A1 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A1 (.I(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__I (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A1 (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__I (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__I (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__I (.I(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A1 (.I(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__I (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A1 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__I (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__I (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A1 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__I (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__I (.I(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__I (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__I (.I(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__I (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__I (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__I (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__I (.I(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A2 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__I (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A2 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A2 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A2 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__A1 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__I (.I(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__I (.I(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A1 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__A1 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A1 (.I(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A1 (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__I (.I(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__I (.I(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A1 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__I (.I(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__I (.I(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__I (.I(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I (.I(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A2 (.I(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A2 (.I(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11297__A2 (.I(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A2 (.I(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A2 (.I(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A2 (.I(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A2 (.I(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A2 (.I(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A1 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__I (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__I (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A1 (.I(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A1 (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__I (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__I (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__I (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__I (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__I (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__I (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A2 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A2 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A2 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__A2 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__I (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__I (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A1 (.I(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__A1 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A1 (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__I (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__I (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A1 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__A1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__I (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__I (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A1 (.I(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__I (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__I (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A2 (.I(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A2 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A2 (.I(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A2 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A2 (.I(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A2 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A2 (.I(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A2 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__CLK (.I(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__CLK (.I(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__CLK (.I(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__CLK (.I(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__CLK (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__CLK (.I(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__CLK (.I(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__CLK (.I(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__CLK (.I(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__CLK (.I(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__CLK (.I(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__CLK (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__CLK (.I(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__CLK (.I(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__CLK (.I(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__CLK (.I(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__CLK (.I(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__CLK (.I(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__D (.I(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__CLK (.I(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__CLK (.I(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__CLK (.I(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__CLK (.I(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__CLK (.I(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__CLK (.I(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__CLK (.I(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__CLK (.I(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__CLK (.I(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__CLK (.I(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__CLK (.I(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__CLK (.I(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__CLK (.I(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__CLK (.I(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__CLK (.I(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__CLK (.I(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__CLK (.I(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__D (.I(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__CLK (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__CLK (.I(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__CLK (.I(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__CLK (.I(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__CLK (.I(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11500__CLK (.I(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__D (.I(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__D (.I(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__D (.I(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11599__D (.I(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__D (.I(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__D (.I(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__D (.I(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__D (.I(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__D (.I(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__CLK (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11639__D (.I(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__D (.I(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__CLK (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__CLK (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__CLK (.I(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11736__CLK (.I(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__CLK (.I(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11792__CLK (.I(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__CLK (.I(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11795__CLK (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11799__CLK (.I(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11823__CLK (.I(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11836__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11881__CLK (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11888__CLK (.I(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11925__CLK (.I(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__CLK (.I(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__CLK (.I(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__CLK (.I(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__CLK (.I(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11974__CLK (.I(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12023__I (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12024__I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12025__I (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12026__I (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__I (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12028__I (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__I (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12030__I (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_137_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_142_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout307_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout308_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold100_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold101_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold102_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold103_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold104_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold105_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold106_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold107_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold108_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold109_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold110_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold111_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold112_I (.I(wbs_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold113_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold114_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold115_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold116_I (.I(wbs_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold117_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold118_I (.I(wbs_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold119_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold120_I (.I(wbs_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold121_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold122_I (.I(wbs_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold123_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold124_I (.I(wbs_adr_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold125_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold126_I (.I(wbs_adr_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold128_I (.I(wbs_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold129_I (.I(wbs_adr_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold130_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold35_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold43_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold50_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold79_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold89_I (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold92_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold93_I (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold94_I (.I(wbs_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold95_I (.I(wbs_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold96_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold97_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold98_I (.I(wbs_adr_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold99_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(bus_in_serial_ports[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(bus_in_serial_ports[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(bus_in_serial_ports[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(bus_in_serial_ports[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(bus_in_serial_ports[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(bus_in_serial_ports[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(bus_in_serial_ports[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(bus_in_sid[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(bus_in_sid[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(bus_in_sid[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(bus_in_gpios[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(bus_in_sid[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(bus_in_sid[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(bus_in_sid[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(bus_in_sid[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(bus_in_sid[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(bus_in_timers[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(bus_in_timers[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(bus_in_timers[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(bus_in_timers[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(bus_in_timers[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(bus_in_gpios[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(bus_in_timers[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(bus_in_timers[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(bus_in_timers[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(bus_in_gpios[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(irqs[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(irqs[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(irqs[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(irqs[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(irqs[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(irqs[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(irqs[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(bus_in_gpios[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(ram_bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(ram_bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(ram_bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(ram_bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(ram_bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(ram_bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(ram_bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(ram_bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(rom_bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(rom_bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(bus_in_gpios[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(rom_bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(rom_bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(rom_bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(rom_bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(rom_bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(rom_bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(bus_in_gpios[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_in_gpios[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(bus_in_gpios[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(bus_in_serial_ports[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap309_I (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output132_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output133_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output134_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output140_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output141_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output142_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output199_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output200_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output209_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output210_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output211_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output212_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output213_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output214_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output215_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output216_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output217_I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output218_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output219_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output220_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output221_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output222_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output223_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output224_I (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output225_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output226_I (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output227_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output228_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output229_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output230_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output231_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output232_I (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output233_I (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output234_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output235_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output236_I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output237_I (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output238_I (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output239_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output240_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output241_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output242_I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output243_I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output244_I (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output245_I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output246_I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output247_I (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output248_I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output249_I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output250_I (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output251_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output252_I (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output253_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output254_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output255_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output256_I (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output266_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output277_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output285_I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output286_I (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output287_I (.I(net287));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output288_I (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output289_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output290_I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output291_I (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output292_I (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output293_I (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer2_I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer5_I (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire298_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire299_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire300_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire301_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire302_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire303_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire304_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire305_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Left_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Left_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Left_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Left_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Left_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Left_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Left_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Left_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Left_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Left_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Left_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Left_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Left_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_668 ();
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _05658_ (.I(\as2650.indirect_cyc ),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05659_ (.I(\as2650.extend ),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05660_ (.A1(_00588_),
    .A2(_00589_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05661_ (.A1(\as2650.instruction_args_latch[13] ),
    .A2(_00590_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05662_ (.I(\as2650.page_reg[0] ),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05663_ (.I(\as2650.indirect_cyc ),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05664_ (.A1(_00593_),
    .A2(\as2650.extend ),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05665_ (.I(\as2650.cycle[9] ),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05666_ (.I(_00595_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05667_ (.I(_00596_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05668_ (.I(_00597_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05669_ (.I(_00598_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05670_ (.A1(_00592_),
    .A2(_00594_),
    .B(_00599_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05671_ (.I(\as2650.relative_cyc ),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05672_ (.I(_00601_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05673_ (.A1(_00602_),
    .A2(_00588_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05674_ (.I(_00603_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05675_ (.I(_00604_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05676_ (.I(_00605_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05677_ (.I(_00606_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _05678_ (.A1(\as2650.relative_cyc ),
    .A2(\as2650.indirect_cyc ),
    .A3(\as2650.cycle[9] ),
    .A4(\as2650.is_interrupt_cycle ),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05679_ (.I(\as2650.cycle[0] ),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05680_ (.A1(_00609_),
    .A2(\as2650.cycle[4] ),
    .A3(\as2650.cycle[6] ),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05681_ (.A1(_00610_),
    .A2(_00608_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05682_ (.I(_00611_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05683_ (.I(_00612_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05684_ (.I(_00613_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05685_ (.I(_00614_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05686_ (.A1(\as2650.indirect_target[13] ),
    .A2(_00607_),
    .B1(_00615_),
    .B2(\as2650.page_reg[0] ),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05687_ (.A1(\as2650.indirect_target[12] ),
    .A2(_00607_),
    .B1(_00615_),
    .B2(\as2650.PC[12] ),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05688_ (.I(_00617_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05689_ (.A1(\as2650.indirect_target[11] ),
    .A2(_00606_),
    .B1(_00614_),
    .B2(\as2650.PC[11] ),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05690_ (.A1(\as2650.indirect_target[10] ),
    .A2(_00606_),
    .B1(_00614_),
    .B2(\as2650.PC[10] ),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05691_ (.A1(\as2650.indirect_target[8] ),
    .A2(_00605_),
    .B1(_00613_),
    .B2(\as2650.PC[8] ),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05692_ (.A1(\as2650.indirect_target[7] ),
    .A2(_00605_),
    .B1(_00613_),
    .B2(\as2650.PC[7] ),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05693_ (.I(\as2650.indirect_target[6] ),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05694_ (.A1(_00601_),
    .A2(_00593_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05695_ (.A1(\as2650.PC[6] ),
    .A2(_00613_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05696_ (.A1(_00623_),
    .A2(_00624_),
    .B(_00625_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05697_ (.A1(\as2650.indirect_target[5] ),
    .A2(_00605_),
    .B1(_00612_),
    .B2(\as2650.PC[5] ),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05698_ (.A1(\as2650.indirect_target[4] ),
    .A2(_00604_),
    .B1(_00612_),
    .B2(\as2650.PC[4] ),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05699_ (.I(\as2650.indirect_target[3] ),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05700_ (.I(_00608_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05701_ (.A1(_00630_),
    .A2(_00610_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05702_ (.I(\as2650.PC[3] ),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _05703_ (.A1(_00629_),
    .A2(_00624_),
    .B1(_00631_),
    .B2(_00632_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05704_ (.A1(\as2650.indirect_target[1] ),
    .A2(_00603_),
    .B1(_00611_),
    .B2(\as2650.PC[1] ),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05705_ (.I(\as2650.cycle[4] ),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05706_ (.I(\as2650.indirect_target[0] ),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05707_ (.A1(_00635_),
    .A2(_00636_),
    .A3(_00604_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05708_ (.A1(\as2650.indirect_target[2] ),
    .A2(_00604_),
    .B1(_00612_),
    .B2(\as2650.PC[2] ),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05709_ (.A1(_00634_),
    .A2(_00637_),
    .A3(_00638_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05710_ (.A1(_00639_),
    .A2(_00633_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05711_ (.A1(_00627_),
    .A2(_00628_),
    .A3(_00640_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05712_ (.A1(_00626_),
    .A2(_00641_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05713_ (.A1(_00621_),
    .A2(_00622_),
    .A3(_00642_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05714_ (.I(_00643_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05715_ (.I(_00644_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05716_ (.A1(\as2650.indirect_target[9] ),
    .A2(_00606_),
    .B1(_00614_),
    .B2(\as2650.PC[9] ),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05717_ (.A1(_00619_),
    .A2(_00620_),
    .A3(_00645_),
    .A4(_00646_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05718_ (.A1(_00618_),
    .A2(_00647_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05719_ (.A1(_00616_),
    .A2(_00648_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05720_ (.I(_00599_),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05721_ (.A1(_00591_),
    .A2(_00600_),
    .B1(_00649_),
    .B2(_00650_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05722_ (.I(_00597_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05723_ (.A1(\as2650.indexed_cyc[1] ),
    .A2(\as2650.indexed_cyc[0] ),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05724_ (.I(_00653_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05725_ (.A1(_00595_),
    .A2(_00654_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05726_ (.I(_00655_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05727_ (.I(_00656_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05728_ (.I(_00657_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05729_ (.I(\as2650.cycle[0] ),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05730_ (.I(_00659_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05731_ (.A1(\as2650.wb_hidden_rom_enable ),
    .A2(\as2650.cpu_hidden_rom_enable ),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05732_ (.I(_00661_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _05733_ (.I(net239),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _05734_ (.A1(net227),
    .A2(net226),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _05735_ (.A1(net225),
    .A2(net224),
    .A3(net223),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05736_ (.A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05737_ (.I0(net39),
    .I1(net51),
    .S(_00666_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05738_ (.A1(net59),
    .A2(_00661_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05739_ (.A1(_00662_),
    .A2(_00667_),
    .B(_00668_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05740_ (.A1(\as2650.insin[1] ),
    .A2(_00659_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05741_ (.A1(_00660_),
    .A2(_00669_),
    .B(_00670_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05742_ (.I(_00671_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05743_ (.I(_00672_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05744_ (.I(_00673_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05745_ (.I(net38),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05746_ (.A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .B(_00675_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05747_ (.A1(_00663_),
    .A2(net50),
    .A3(_00664_),
    .A4(_00665_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05748_ (.A1(_00676_),
    .A2(_00677_),
    .B(_00662_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05749_ (.A1(net58),
    .A2(_00661_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05750_ (.A1(\as2650.insin[0] ),
    .A2(_00659_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05751_ (.A1(_00659_),
    .A2(_00678_),
    .A3(_00679_),
    .B(_00680_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05752_ (.I(_00681_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05753_ (.I(_00682_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05754_ (.I(_00683_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05755_ (.I(\as2650.debug_psl[4] ),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05756_ (.I(_00685_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05757_ (.I(_00686_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05758_ (.I(_00687_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05759_ (.I(\as2650.debug_psl[4] ),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05760_ (.I(_00689_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05761_ (.I(_00690_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05762_ (.A1(_00691_),
    .A2(\as2650.regs[0][7] ),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05763_ (.A1(_00688_),
    .A2(\as2650.regs[4][7] ),
    .B(_00692_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05764_ (.I(_00693_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05765_ (.I(_00694_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05766_ (.I(\as2650.debug_psl[4] ),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05767_ (.I0(\as2650.regs[1][7] ),
    .I1(\as2650.regs[5][7] ),
    .S(_00696_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05768_ (.I(_00697_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _05769_ (.I(_00698_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05770_ (.A1(_00684_),
    .A2(_00699_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05771_ (.A1(_00684_),
    .A2(_00695_),
    .B(_00700_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05772_ (.I(_00673_),
    .Z(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05773_ (.I(\as2650.regs[2][7] ),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05774_ (.A1(_00688_),
    .A2(\as2650.regs[6][7] ),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05775_ (.A1(_00688_),
    .A2(_00703_),
    .B(_00704_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05776_ (.I(_00705_),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05777_ (.I(_00687_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05778_ (.I(_00706_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05779_ (.I(\as2650.regs[3][7] ),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05780_ (.A1(_00707_),
    .A2(\as2650.regs[7][7] ),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05781_ (.A1(_00707_),
    .A2(_00708_),
    .B(_00709_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05782_ (.I(_00681_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05783_ (.I(_00711_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05784_ (.I0(net203),
    .I1(_00710_),
    .S(_00712_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05785_ (.A1(_00702_),
    .A2(_00713_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05786_ (.A1(_00674_),
    .A2(_00701_),
    .B(_00714_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05787_ (.I(_00715_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05788_ (.A1(_00622_),
    .A2(_00642_),
    .B(_00598_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05789_ (.A1(_00622_),
    .A2(_00642_),
    .B(_00717_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _05790_ (.A1(_00652_),
    .A2(\as2650.instruction_args_latch[7] ),
    .B1(_00658_),
    .B2(_00716_),
    .C(_00718_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05791_ (.I(_00719_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05792_ (.I(\as2650.cycle[9] ),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05793_ (.I(\as2650.debug_psl[4] ),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05794_ (.I(_00722_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05795_ (.I(\as2650.regs[0][0] ),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05796_ (.A1(_00685_),
    .A2(_00724_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05797_ (.A1(_00723_),
    .A2(\as2650.regs[4][0] ),
    .B(_00725_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05798_ (.I(_00726_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05799_ (.I(_00722_),
    .Z(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05800_ (.I0(\as2650.regs[1][0] ),
    .I1(\as2650.regs[5][0] ),
    .S(_00728_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05801_ (.I(net353),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05802_ (.I0(_00727_),
    .I1(_00729_),
    .S(_00730_),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05803_ (.A1(_00689_),
    .A2(\as2650.regs[2][0] ),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05804_ (.I(_00722_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05805_ (.A1(_00733_),
    .A2(\as2650.regs[6][0] ),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05806_ (.A1(_00732_),
    .A2(_00734_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05807_ (.I(_00735_),
    .ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _05808_ (.I(_00723_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05809_ (.I(\as2650.regs[3][0] ),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05810_ (.A1(_00728_),
    .A2(\as2650.regs[7][0] ),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05811_ (.A1(_00736_),
    .A2(_00737_),
    .B(_00738_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05812_ (.I0(net195),
    .I1(_00739_),
    .S(_00730_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05813_ (.I0(_00731_),
    .I1(_00740_),
    .S(_00671_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _05814_ (.A1(\as2650.instruction_args_latch[0] ),
    .A2(_00721_),
    .A3(_00654_),
    .A4(_00741_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05815_ (.A1(_00595_),
    .A2(_00653_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05816_ (.I(_00743_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05817_ (.I(\as2650.regs[0][1] ),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05818_ (.A1(_00685_),
    .A2(_00745_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05819_ (.A1(_00696_),
    .A2(\as2650.regs[4][1] ),
    .B(_00746_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05820_ (.I0(\as2650.regs[1][1] ),
    .I1(\as2650.regs[5][1] ),
    .S(_00722_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _05821_ (.I(_00748_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05822_ (.I0(_00747_),
    .I1(_00749_),
    .S(_00730_),
    .Z(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05823_ (.A1(_00690_),
    .A2(\as2650.regs[2][1] ),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05824_ (.A1(_00696_),
    .A2(\as2650.regs[6][1] ),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05825_ (.A1(_00751_),
    .A2(_00752_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05826_ (.I(\as2650.regs[3][1] ),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05827_ (.A1(_00733_),
    .A2(\as2650.regs[7][1] ),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05828_ (.A1(_00696_),
    .A2(_00754_),
    .B(_00755_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05829_ (.I(_00756_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05830_ (.I0(_00753_),
    .I1(_00757_),
    .S(_00730_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05831_ (.I0(_00750_),
    .I1(_00758_),
    .S(_00671_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05832_ (.I(_00759_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05833_ (.A1(_00635_),
    .A2(\as2650.indirect_target[0] ),
    .A3(_00603_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05834_ (.A1(_00634_),
    .A2(_00761_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05835_ (.A1(\as2650.cycle[9] ),
    .A2(\as2650.instruction_args_latch[1] ),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05836_ (.A1(_00595_),
    .A2(_00762_),
    .B(_00763_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05837_ (.I(_00764_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05838_ (.A1(_00744_),
    .A2(_00760_),
    .B(_00765_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05839_ (.A1(_00743_),
    .A2(_00759_),
    .A3(_00765_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05840_ (.A1(_00742_),
    .A2(_00766_),
    .B(_00767_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05841_ (.A1(_00689_),
    .A2(\as2650.regs[0][2] ),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05842_ (.A1(_00686_),
    .A2(\as2650.regs[4][2] ),
    .B(_00769_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05843_ (.I0(\as2650.regs[1][2] ),
    .I1(\as2650.regs[5][2] ),
    .S(_00736_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _05844_ (.I(_00771_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05845_ (.I0(_00770_),
    .I1(_00772_),
    .S(_00711_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05846_ (.A1(_00690_),
    .A2(\as2650.regs[2][2] ),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05847_ (.I(_00733_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05848_ (.A1(_00775_),
    .A2(\as2650.regs[6][2] ),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05849_ (.A1(_00774_),
    .A2(_00776_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05850_ (.I(_00777_),
    .ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05851_ (.I(_00733_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05852_ (.I(\as2650.regs[3][2] ),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05853_ (.A1(_00728_),
    .A2(\as2650.regs[7][2] ),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05854_ (.A1(_00778_),
    .A2(_00779_),
    .B(_00780_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05855_ (.I(_00781_),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05856_ (.I(net206),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05857_ (.A1(_00711_),
    .A2(_00782_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05858_ (.A1(_00683_),
    .A2(net197),
    .B(_00783_),
    .C(_00672_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05859_ (.A1(_00673_),
    .A2(_00773_),
    .B(_00784_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05860_ (.A1(_00634_),
    .A2(_00637_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05861_ (.A1(_00786_),
    .A2(_00638_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05862_ (.A1(_00721_),
    .A2(\as2650.instruction_args_latch[2] ),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05863_ (.A1(_00596_),
    .A2(_00787_),
    .B(_00788_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05864_ (.A1(_00656_),
    .A2(_00785_),
    .B(_00789_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05865_ (.A1(_00655_),
    .A2(_00785_),
    .A3(_00789_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05866_ (.A1(_00768_),
    .A2(_00790_),
    .B(_00791_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05867_ (.I0(\as2650.regs[0][3] ),
    .I1(\as2650.regs[4][3] ),
    .S(_00685_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05868_ (.I(_00793_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05869_ (.I0(\as2650.regs[1][3] ),
    .I1(\as2650.regs[5][3] ),
    .S(_00723_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _05870_ (.I(_00795_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05871_ (.I0(_00794_),
    .I1(_00796_),
    .S(_00682_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05872_ (.A1(_00690_),
    .A2(\as2650.regs[2][3] ),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05873_ (.A1(_00778_),
    .A2(\as2650.regs[6][3] ),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _05874_ (.A1(_00798_),
    .A2(_00799_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05875_ (.I(\as2650.regs[3][3] ),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05876_ (.A1(_00728_),
    .A2(\as2650.regs[7][3] ),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05877_ (.A1(_00778_),
    .A2(_00801_),
    .B(_00802_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05878_ (.I(_00803_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05879_ (.I0(_00800_),
    .I1(_00804_),
    .S(_00682_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05880_ (.I0(_00797_),
    .I1(_00805_),
    .S(_00672_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05881_ (.A1(_00743_),
    .A2(_00806_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _05882_ (.A1(_00633_),
    .A2(_00639_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05883_ (.A1(_00721_),
    .A2(\as2650.instruction_args_latch[3] ),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05884_ (.A1(_00721_),
    .A2(_00808_),
    .B(_00809_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05885_ (.A1(_00807_),
    .A2(_00810_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05886_ (.A1(_00807_),
    .A2(_00810_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05887_ (.A1(_00792_),
    .A2(_00811_),
    .B(_00812_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05888_ (.I(\as2650.regs[0][4] ),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05889_ (.A1(_00686_),
    .A2(_00814_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05890_ (.A1(_00736_),
    .A2(\as2650.regs[4][4] ),
    .B(_00815_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05891_ (.I(_00816_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05892_ (.I(_00817_),
    .Z(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05893_ (.I(_00818_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05894_ (.I0(\as2650.regs[1][4] ),
    .I1(\as2650.regs[5][4] ),
    .S(_00775_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05895_ (.I(_00820_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _05896_ (.I(_00821_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05897_ (.A1(_00712_),
    .A2(_00822_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05898_ (.A1(_00712_),
    .A2(_00819_),
    .B(_00823_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05899_ (.I(\as2650.regs[2][4] ),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05900_ (.I(_00775_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05901_ (.A1(_00826_),
    .A2(\as2650.regs[6][4] ),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05902_ (.A1(_00688_),
    .A2(_00825_),
    .B(_00827_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05903_ (.I(_00828_),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05904_ (.I(\as2650.regs[3][4] ),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05905_ (.A1(_00826_),
    .A2(\as2650.regs[7][4] ),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05906_ (.A1(_00706_),
    .A2(_00829_),
    .B(_00830_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05907_ (.I(_00831_),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05908_ (.I(_00682_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05909_ (.I0(net200),
    .I1(net208),
    .S(_00832_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05910_ (.A1(_00702_),
    .A2(_00833_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05911_ (.A1(_00702_),
    .A2(_00824_),
    .B(_00834_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05912_ (.I(_00596_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05913_ (.A1(_00628_),
    .A2(_00640_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05914_ (.A1(_00836_),
    .A2(\as2650.instruction_args_latch[4] ),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05915_ (.A1(_00836_),
    .A2(_00837_),
    .B(_00838_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05916_ (.A1(_00657_),
    .A2(_00835_),
    .B(_00839_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05917_ (.A1(_00657_),
    .A2(_00835_),
    .A3(_00839_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05918_ (.A1(_00813_),
    .A2(_00840_),
    .B(_00841_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05919_ (.I(_00686_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05920_ (.I(\as2650.regs[2][5] ),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05921_ (.A1(_00687_),
    .A2(\as2650.regs[6][5] ),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05922_ (.A1(_00843_),
    .A2(_00844_),
    .B(_00845_),
    .ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05923_ (.I(net201),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05924_ (.I(\as2650.regs[3][5] ),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05925_ (.A1(_00843_),
    .A2(\as2650.regs[7][5] ),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05926_ (.A1(_00826_),
    .A2(_00847_),
    .B(_00848_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05927_ (.A1(_00711_),
    .A2(_00849_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05928_ (.A1(_00832_),
    .A2(_00846_),
    .B(_00850_),
    .C(_00672_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05929_ (.I(\as2650.regs[0][5] ),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05930_ (.A1(_00778_),
    .A2(_00852_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05931_ (.A1(_00775_),
    .A2(\as2650.regs[4][5] ),
    .B(_00853_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05932_ (.I(_00854_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05933_ (.I0(\as2650.regs[1][5] ),
    .I1(\as2650.regs[5][5] ),
    .S(_00736_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05934_ (.I(_00856_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05935_ (.A1(_00683_),
    .A2(_00857_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05936_ (.I(_00661_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05937_ (.I0(net59),
    .I1(_00667_),
    .S(_00859_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05938_ (.A1(_00609_),
    .A2(_00860_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05939_ (.A1(_00670_),
    .A2(_00861_),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05940_ (.A1(_00832_),
    .A2(_00855_),
    .B(_00858_),
    .C(_00862_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05941_ (.A1(_00851_),
    .A2(_00863_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05942_ (.A1(_00656_),
    .A2(_00864_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05943_ (.A1(_00628_),
    .A2(_00640_),
    .B(_00627_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05944_ (.A1(_00596_),
    .A2(_00641_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05945_ (.A1(_00836_),
    .A2(\as2650.instruction_args_latch[5] ),
    .B1(_00866_),
    .B2(_00867_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05946_ (.A1(_00865_),
    .A2(_00868_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05947_ (.A1(_00865_),
    .A2(_00868_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05948_ (.A1(_00842_),
    .A2(_00869_),
    .B(_00870_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05949_ (.I(\as2650.regs[0][6] ),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05950_ (.A1(_00687_),
    .A2(_00872_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05951_ (.A1(_00843_),
    .A2(\as2650.regs[4][6] ),
    .B(_00873_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05952_ (.I(_00874_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05953_ (.I(_00875_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05954_ (.I0(\as2650.regs[1][6] ),
    .I1(\as2650.regs[5][6] ),
    .S(_00723_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05955_ (.I(_00877_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05956_ (.I(_00878_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05957_ (.A1(_00832_),
    .A2(_00879_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05958_ (.A1(_00712_),
    .A2(_00876_),
    .B(_00880_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05959_ (.I(\as2650.regs[2][6] ),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05960_ (.A1(_00826_),
    .A2(\as2650.regs[6][6] ),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05961_ (.A1(_00706_),
    .A2(_00882_),
    .B(_00883_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05962_ (.I(_00884_),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05963_ (.I(\as2650.regs[3][6] ),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05964_ (.A1(_00843_),
    .A2(\as2650.regs[7][6] ),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05965_ (.A1(_00706_),
    .A2(_00885_),
    .B(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05966_ (.I(_00887_),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05967_ (.I0(net202),
    .I1(net211),
    .S(_00683_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05968_ (.A1(_00673_),
    .A2(_00888_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05969_ (.A1(_00702_),
    .A2(_00881_),
    .B(_00889_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05970_ (.A1(_00656_),
    .A2(_00890_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05971_ (.A1(_00626_),
    .A2(_00641_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05972_ (.A1(_00836_),
    .A2(\as2650.instruction_args_latch[6] ),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05973_ (.A1(_00597_),
    .A2(_00892_),
    .B(_00893_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05974_ (.A1(_00891_),
    .A2(_00894_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05975_ (.A1(_00652_),
    .A2(\as2650.instruction_args_latch[7] ),
    .A3(_00654_),
    .A4(_00715_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05976_ (.A1(_00657_),
    .A2(_00890_),
    .A3(_00894_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _05977_ (.A1(_00871_),
    .A2(_00895_),
    .B(_00896_),
    .C(_00897_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _05978_ (.I(\as2650.instruction_args_latch[8] ),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05979_ (.A1(_00599_),
    .A2(_00899_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05980_ (.A1(_00622_),
    .A2(_00642_),
    .B(_00621_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05981_ (.A1(_00599_),
    .A2(_00645_),
    .A3(_00901_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05982_ (.A1(_00900_),
    .A2(_00902_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05983_ (.I(_00597_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05984_ (.A1(_00645_),
    .A2(_00646_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05985_ (.A1(_00644_),
    .A2(_00646_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05986_ (.A1(_00652_),
    .A2(_00906_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05987_ (.A1(_00904_),
    .A2(\as2650.instruction_args_latch[9] ),
    .B1(_00905_),
    .B2(_00907_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05988_ (.I(_00908_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05989_ (.A1(_00720_),
    .A2(_00898_),
    .A3(_00903_),
    .A4(_00909_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05990_ (.I(_00652_),
    .Z(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05991_ (.A1(_00620_),
    .A2(_00906_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05992_ (.A1(_00904_),
    .A2(_00912_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05993_ (.A1(_00911_),
    .A2(\as2650.instruction_args_latch[10] ),
    .B(_00913_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05994_ (.I(_00904_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05995_ (.A1(_00620_),
    .A2(_00645_),
    .A3(_00646_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05996_ (.A1(_00619_),
    .A2(_00916_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05997_ (.A1(_00911_),
    .A2(_00917_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05998_ (.A1(_00915_),
    .A2(\as2650.instruction_args_latch[11] ),
    .B(_00918_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05999_ (.A1(_00618_),
    .A2(_00647_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06000_ (.A1(_00911_),
    .A2(_00648_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06001_ (.A1(_00915_),
    .A2(\as2650.instruction_args_latch[12] ),
    .B1(_00920_),
    .B2(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06002_ (.A1(_00910_),
    .A2(_00914_),
    .A3(_00919_),
    .A4(_00922_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06003_ (.I(_00915_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06004_ (.I(\as2650.instruction_args_latch[14] ),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06005_ (.A1(_00925_),
    .A2(_00594_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06006_ (.A1(\as2650.page_reg[1] ),
    .A2(_00594_),
    .B(_00926_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06007_ (.A1(_00618_),
    .A2(_00647_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06008_ (.A1(_00616_),
    .A2(_00928_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06009_ (.I(\as2650.indirect_target[14] ),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06010_ (.I(_00631_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06011_ (.I(\as2650.page_reg[1] ),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06012_ (.A1(_00930_),
    .A2(_00624_),
    .B1(_00931_),
    .B2(_00932_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06013_ (.A1(_00929_),
    .A2(_00933_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06014_ (.A1(_00924_),
    .A2(_00934_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06015_ (.A1(_00924_),
    .A2(_00927_),
    .B(_00935_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06016_ (.A1(_00651_),
    .A2(_00923_),
    .A3(_00936_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06017_ (.I(_00924_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06018_ (.I(\as2650.instruction_args_latch[15] ),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06019_ (.I(_00594_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06020_ (.A1(\as2650.page_reg[2] ),
    .A2(_00940_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06021_ (.A1(_00939_),
    .A2(_00940_),
    .B(_00941_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06022_ (.A1(_00929_),
    .A2(_00933_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06023_ (.I(_00615_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06024_ (.A1(\as2650.indirect_target[15] ),
    .A2(_00607_),
    .B1(_00944_),
    .B2(\as2650.page_reg[2] ),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06025_ (.A1(_00943_),
    .A2(_00945_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06026_ (.A1(_00943_),
    .A2(_00945_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06027_ (.A1(_00924_),
    .A2(_00947_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06028_ (.A1(_00938_),
    .A2(_00942_),
    .B1(_00946_),
    .B2(_00948_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06029_ (.A1(_00937_),
    .A2(_00949_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06030_ (.I(_00950_),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06031_ (.I(net225),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06032_ (.A1(_00651_),
    .A2(_00923_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06033_ (.I(_00952_),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06034_ (.I(_00910_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06035_ (.I(_00914_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06036_ (.A1(net222),
    .A2(_00953_),
    .A3(_00954_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06037_ (.I(net236),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06038_ (.A1(_00720_),
    .A2(_00898_),
    .A3(_00903_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06039_ (.A1(_00956_),
    .A2(_00957_),
    .A3(_00908_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06040_ (.A1(_00720_),
    .A2(_00898_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06041_ (.A1(net235),
    .A2(_00959_),
    .A3(_00903_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06042_ (.A1(_00955_),
    .A2(_00958_),
    .A3(_00960_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06043_ (.A1(_00953_),
    .A2(_00954_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06044_ (.A1(net223),
    .A2(_00962_),
    .A3(_00919_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06045_ (.A1(_00951_),
    .A2(net244),
    .B(_00961_),
    .C(_00963_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06046_ (.A1(_00651_),
    .A2(_00923_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06047_ (.A1(_00651_),
    .A2(_00923_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06048_ (.A1(_00953_),
    .A2(_00954_),
    .A3(_00919_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06049_ (.A1(net224),
    .A2(_00967_),
    .A3(_00922_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06050_ (.A1(net225),
    .A2(_00965_),
    .A3(_00966_),
    .B(_00968_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06051_ (.A1(net226),
    .A2(_00965_),
    .A3(_00936_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06052_ (.I(net227),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06053_ (.A1(_00971_),
    .A2(_00937_),
    .A3(_00949_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _06054_ (.A1(_00964_),
    .A2(_00969_),
    .A3(_00970_),
    .A4(_00972_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06055_ (.I(_00973_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06056_ (.I(_00974_),
    .Z(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06057_ (.I(_00975_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06058_ (.I(\as2650.cycle[8] ),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06059_ (.I(_00609_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06060_ (.I(_00978_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06061_ (.I(_00979_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06062_ (.I(_00635_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06063_ (.I(_00981_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06064_ (.I(\as2650.cycle[6] ),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06065_ (.A1(_00980_),
    .A2(_00982_),
    .A3(_00983_),
    .A4(_00630_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06066_ (.A1(\as2650.cycle[2] ),
    .A2(_00977_),
    .A3(_00984_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06067_ (.A1(_00976_),
    .A2(_00985_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06068_ (.I(_00986_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06069_ (.I(_00987_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06070_ (.I(_00988_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06071_ (.I(_00989_),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06072_ (.A1(_00965_),
    .A2(_00936_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06073_ (.I(_00990_),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06074_ (.A1(_00967_),
    .A2(_00922_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06075_ (.I(_00991_),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06076_ (.A1(_00962_),
    .A2(_00919_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06077_ (.I(_00992_),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06078_ (.A1(_00953_),
    .A2(_00954_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06079_ (.I(_00993_),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06080_ (.A1(_00957_),
    .A2(_00908_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06081_ (.I(_00994_),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06082_ (.A1(_00959_),
    .A2(_00903_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06083_ (.I(_00995_),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06084_ (.I(_00698_),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06085_ (.I(_00996_),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06086_ (.I(_00878_),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06087_ (.I(_00857_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06088_ (.I(_00997_),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06089_ (.I(_00821_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06090_ (.I(_00998_),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06091_ (.I(_00795_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06092_ (.I(_00999_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06093_ (.I(_01000_),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06094_ (.I(_00771_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06095_ (.I(_01001_),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06096_ (.I(_00748_),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06097_ (.I(_01002_),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06098_ (.I(_01003_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06099_ (.I(_01004_),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06100_ (.I(_00729_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06101_ (.I(_01005_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06102_ (.I(_01006_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06103_ (.I(_01007_),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06104_ (.I(_00695_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06105_ (.I(_01008_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06106_ (.I(_01009_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06107_ (.I(_01010_),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06108_ (.I(_00876_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06109_ (.I(_01011_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06110_ (.I(_01012_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06111_ (.I(_01013_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06112_ (.I(_01014_),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06113_ (.I(_00854_),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06114_ (.I(_01015_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06115_ (.I(_01016_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06116_ (.I(_01017_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06117_ (.I(_01018_),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06118_ (.I(_00819_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06119_ (.I(_01019_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06120_ (.I(_01020_),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06121_ (.A1(wb_reset_override),
    .A2(wb_reset_override_en),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06122_ (.A1(wb_reset_override_en),
    .A2(net33),
    .B(_01021_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06123_ (.A1(net66),
    .A2(_01022_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06124_ (.I(_01023_),
    .ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06125_ (.A1(_00871_),
    .A2(_00895_),
    .B(_00897_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06126_ (.A1(_00720_),
    .A2(_00896_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06127_ (.A1(_01024_),
    .A2(_01025_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06128_ (.I(_01026_),
    .ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06129_ (.I(net229),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06130_ (.I(_00658_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06131_ (.A1(_01028_),
    .A2(_00785_),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06132_ (.A1(_01029_),
    .A2(_00789_),
    .A3(_00768_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06133_ (.I(_01030_),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06134_ (.A1(_00674_),
    .A2(_00758_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06135_ (.A1(_00862_),
    .A2(_00750_),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06136_ (.A1(_01031_),
    .A2(_01032_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06137_ (.A1(_00658_),
    .A2(_01033_),
    .A3(_00764_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06138_ (.I(\as2650.instruction_args_latch[0] ),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06139_ (.A1(_01035_),
    .A2(_00911_),
    .A3(_00654_),
    .A4(_00741_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06140_ (.A1(_01034_),
    .A2(_01036_),
    .A3(_00766_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06141_ (.A1(_00658_),
    .A2(_01033_),
    .B(_00764_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06142_ (.A1(_00767_),
    .A2(_01038_),
    .B(_00742_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06143_ (.A1(_01037_),
    .A2(_01039_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06144_ (.I(_01040_),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06145_ (.A1(net228),
    .A2(net247),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06146_ (.A1(\as2650.PC[0] ),
    .A2(_00615_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06147_ (.A1(_00636_),
    .A2(_00607_),
    .B1(_00630_),
    .B2(_00635_),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06148_ (.A1(_01042_),
    .A2(_01043_),
    .B(_00904_),
    .C(_00761_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06149_ (.A1(_01035_),
    .A2(_00915_),
    .B1(_01028_),
    .B2(_00741_),
    .C(_01044_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06150_ (.A1(_00742_),
    .A2(_01045_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06151_ (.I(_01046_),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06152_ (.A1(net221),
    .A2(net240),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06153_ (.A1(_01027_),
    .A2(_01030_),
    .B(_01041_),
    .C(_01047_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06154_ (.A1(_00792_),
    .A2(_00811_),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06155_ (.I(_01049_),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06156_ (.A1(net230),
    .A2(net249),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06157_ (.A1(_01027_),
    .A2(net248),
    .B(_01048_),
    .C(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06158_ (.A1(_01028_),
    .A2(_00835_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06159_ (.A1(_01052_),
    .A2(_00839_),
    .A3(_00813_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06160_ (.I(_01053_),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06161_ (.A1(net231),
    .A2(net250),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06162_ (.A1(_01051_),
    .A2(_01054_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06163_ (.A1(net349),
    .A2(_00869_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06164_ (.I(_01056_),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06165_ (.A1(net232),
    .A2(net251),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06166_ (.A1(_00871_),
    .A2(_00895_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06167_ (.I(_01058_),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06168_ (.A1(net233),
    .A2(net252),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06169_ (.A1(net234),
    .A2(_01026_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _06170_ (.A1(_01055_),
    .A2(_01057_),
    .A3(_01059_),
    .A4(_01060_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06171_ (.I(_01061_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06172_ (.I(_01062_),
    .Z(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06173_ (.I(_01063_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06174_ (.A1(_00985_),
    .A2(_01064_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06175_ (.A1(_00976_),
    .A2(_01065_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06176_ (.I(_01066_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06177_ (.I(_01067_),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06178_ (.I(_01068_),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06179_ (.I(_00662_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06180_ (.I(_01069_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06181_ (.I(_01070_),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06182_ (.A1(net48),
    .A2(net47),
    .A3(net49),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06183_ (.A1(net44),
    .A2(net43),
    .A3(net46),
    .A4(net45),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06184_ (.A1(_01071_),
    .A2(_01072_),
    .B(\as2650.debug_psu[5] ),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06185_ (.I(_01073_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _06186_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(net256),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06187_ (.I(_01075_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06188_ (.I(_01076_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06189_ (.I(_01077_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06190_ (.I(_01078_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06191_ (.I(_01079_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06192_ (.I(_01080_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06193_ (.I(\as2650.extend ),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06194_ (.I(_01082_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06195_ (.I(_00862_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06196_ (.I(_01084_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06197_ (.A1(_00678_),
    .A2(_00679_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06198_ (.A1(_00979_),
    .A2(_01086_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06199_ (.A1(_00680_),
    .A2(_01087_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06200_ (.I(_00666_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06201_ (.I0(net41),
    .I1(net53),
    .S(_01089_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _06202_ (.I0(net61),
    .I1(_01090_),
    .S(_00859_),
    .Z(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _06203_ (.I0(\as2650.insin[3] ),
    .I1(_01091_),
    .S(_00609_),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06204_ (.I0(net40),
    .I1(net52),
    .S(_01089_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06205_ (.A1(net60),
    .A2(_00859_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06206_ (.A1(_00662_),
    .A2(_01093_),
    .B(_01094_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06207_ (.A1(\as2650.insin[2] ),
    .A2(_00660_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06208_ (.A1(_00660_),
    .A2(_01095_),
    .B(_01096_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06209_ (.A1(_01092_),
    .A2(_01097_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06210_ (.I(_01098_),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06211_ (.I(_01099_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06212_ (.I(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06213_ (.I(_01101_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06214_ (.A1(_01085_),
    .A2(_01088_),
    .A3(_01102_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06215_ (.I(_01103_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06216_ (.I(_01089_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06217_ (.I(net57),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06218_ (.A1(_01106_),
    .A2(_01105_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06219_ (.A1(net36),
    .A2(_01105_),
    .B(_01107_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06220_ (.A1(net65),
    .A2(_01069_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06221_ (.A1(_01069_),
    .A2(_01108_),
    .B(_01109_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06222_ (.A1(_00978_),
    .A2(_01110_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06223_ (.I(_00660_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06224_ (.A1(\as2650.insin[7] ),
    .A2(_01112_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06225_ (.A1(_01111_),
    .A2(_01113_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06226_ (.I(_01114_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06227_ (.I(_01089_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06228_ (.I(net56),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06229_ (.A1(_01117_),
    .A2(_01105_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06230_ (.A1(net35),
    .A2(_01116_),
    .B(_01118_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06231_ (.A1(net64),
    .A2(_01069_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06232_ (.A1(_01070_),
    .A2(_01119_),
    .B(_01120_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06233_ (.A1(_00978_),
    .A2(_01121_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06234_ (.A1(\as2650.insin[6] ),
    .A2(_01112_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06235_ (.A1(_01122_),
    .A2(_01123_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06236_ (.I(_01124_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06237_ (.A1(_01115_),
    .A2(_01125_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06238_ (.I(_01126_),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06239_ (.I(_01112_),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06240_ (.A1(\as2650.insin[5] ),
    .A2(_01128_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06241_ (.I(net55),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06242_ (.A1(_01130_),
    .A2(_01116_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06243_ (.A1(net34),
    .A2(_01116_),
    .B(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06244_ (.A1(net63),
    .A2(net139),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06245_ (.A1(net139),
    .A2(_01132_),
    .B(_01133_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06246_ (.A1(_00979_),
    .A2(_01134_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06247_ (.A1(_01129_),
    .A2(_01135_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06248_ (.A1(\as2650.insin[4] ),
    .A2(_01112_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06249_ (.I(net54),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06250_ (.A1(_01138_),
    .A2(_01105_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06251_ (.A1(net42),
    .A2(_01116_),
    .B(_01139_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06252_ (.A1(net62),
    .A2(_01070_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06253_ (.A1(_01070_),
    .A2(_01140_),
    .B(_01141_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06254_ (.A1(_00978_),
    .A2(_01142_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06255_ (.A1(_01137_),
    .A2(_01143_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06256_ (.I(_01144_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06257_ (.A1(_01136_),
    .A2(_01145_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06258_ (.A1(_01083_),
    .A2(_01104_),
    .A3(_01127_),
    .A4(_01146_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06259_ (.I(_01147_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06260_ (.A1(_01128_),
    .A2(_00974_),
    .A3(_01062_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06261_ (.I(_01149_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06262_ (.I(_01150_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06263_ (.I(_01151_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06264_ (.A1(_01148_),
    .A2(_01152_),
    .B(\as2650.cycle[11] ),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06265_ (.A1(\as2650.cycle[11] ),
    .A2(_01074_),
    .B(_01081_),
    .C(_01153_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06266_ (.I(_00859_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06267_ (.A1(net61),
    .A2(_01154_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06268_ (.A1(net139),
    .A2(_01090_),
    .B(_01155_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06269_ (.A1(_00979_),
    .A2(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06270_ (.A1(\as2650.insin[3] ),
    .A2(_00980_),
    .B(_01157_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06271_ (.I(_01158_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06272_ (.I(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06273_ (.I(_01097_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06274_ (.A1(_01082_),
    .A2(_01161_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06275_ (.A1(_01160_),
    .A2(_01162_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06276_ (.A1(_00593_),
    .A2(_01163_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06277_ (.I(_00983_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06278_ (.I(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06279_ (.I(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06280_ (.I(_01167_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _06281_ (.A1(_01061_),
    .A2(_00973_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06282_ (.I(_01169_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06283_ (.I(_01170_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06284_ (.I(_01171_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06285_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(net350),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06286_ (.I(_01173_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06287_ (.I(_01174_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06288_ (.I(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06289_ (.I(_01128_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06290_ (.A1(_00973_),
    .A2(_01061_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06291_ (.I(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06292_ (.I(_01179_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06293_ (.I(\as2650.cycle[11] ),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06294_ (.A1(_01177_),
    .A2(_01180_),
    .B(_01181_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06295_ (.A1(_01073_),
    .A2(_01182_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06296_ (.A1(_01176_),
    .A2(_01183_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06297_ (.A1(_01172_),
    .A2(_01184_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06298_ (.I(_01185_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06299_ (.I(_01161_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06300_ (.A1(_01160_),
    .A2(_01187_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06301_ (.A1(_00601_),
    .A2(_01188_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06302_ (.I(_01189_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06303_ (.I(_01190_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06304_ (.A1(_01168_),
    .A2(_01186_),
    .A3(_01191_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06305_ (.I(_00982_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06306_ (.I(_01193_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06307_ (.I(_01180_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06308_ (.I(_01195_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06309_ (.I(_01196_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06310_ (.A1(_01197_),
    .A2(_01184_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06311_ (.A1(_01194_),
    .A2(_01198_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06312_ (.A1(_01164_),
    .A2(_01192_),
    .B(_01199_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06313_ (.I(_01182_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06314_ (.I(_01079_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06315_ (.A1(_01074_),
    .A2(_01200_),
    .B(_01201_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06316_ (.A1(\as2650.cycle[5] ),
    .A2(_01202_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06317_ (.I(_01203_),
    .Z(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06318_ (.I(_00980_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06319_ (.I(_01204_),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06320_ (.I(_01205_),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06321_ (.I(_01206_),
    .Z(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06322_ (.A1(_01129_),
    .A2(_01135_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06323_ (.I(_01208_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06324_ (.A1(_01137_),
    .A2(_01143_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06325_ (.I(_01210_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06326_ (.A1(_01209_),
    .A2(_01211_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06327_ (.I(_01212_),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06328_ (.A1(_01158_),
    .A2(_01162_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06329_ (.I(_01214_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06330_ (.A1(_01213_),
    .A2(_01215_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06331_ (.A1(_01207_),
    .A2(_01186_),
    .A3(_01216_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06332_ (.I(_01217_),
    .Z(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06333_ (.I(_00938_),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06334_ (.I(_01092_),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06335_ (.I(_01211_),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06336_ (.A1(_01219_),
    .A2(_01220_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06337_ (.A1(_00981_),
    .A2(_01221_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06338_ (.A1(_00939_),
    .A2(_00590_),
    .A3(_01159_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06339_ (.I(_01083_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06340_ (.I(_01224_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06341_ (.I(_00674_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06342_ (.I(_01102_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06343_ (.I(_01227_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06344_ (.A1(_01111_),
    .A2(_01113_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06345_ (.I(_01229_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06346_ (.I(_01230_),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06347_ (.A1(_01122_),
    .A2(_01123_),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06348_ (.I(_01232_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06349_ (.A1(_01231_),
    .A2(_01233_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06350_ (.I(_01234_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06351_ (.I(_01136_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06352_ (.I(_01236_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06353_ (.A1(_01237_),
    .A2(_01211_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06354_ (.A1(_01235_),
    .A2(_01238_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06355_ (.I(_01239_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06356_ (.A1(_01225_),
    .A2(_01226_),
    .A3(_01228_),
    .A4(_01240_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06357_ (.A1(_01177_),
    .A2(_01241_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06358_ (.I(_01242_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06359_ (.A1(_01222_),
    .A2(_01223_),
    .B(_01243_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06360_ (.A1(_01218_),
    .A2(_01198_),
    .B1(_01186_),
    .B2(_01244_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06361_ (.I(_01245_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06362_ (.A1(\as2650.cycle[7] ),
    .A2(_01202_),
    .Z(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06363_ (.I(_01246_),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06364_ (.A1(\as2650.cycle[2] ),
    .A2(_01202_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06365_ (.I(_01247_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06366_ (.I(\as2650.cycle[1] ),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06367_ (.A1(_01248_),
    .A2(_01184_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06368_ (.A1(_01185_),
    .A2(_01241_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06369_ (.I(_01163_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06370_ (.I(_01225_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06371_ (.A1(_01159_),
    .A2(_01187_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06372_ (.A1(_01083_),
    .A2(_01252_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06373_ (.I(_01253_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06374_ (.I(_01145_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06375_ (.A1(_01114_),
    .A2(_01232_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06376_ (.A1(_01255_),
    .A2(_01256_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06377_ (.A1(_01219_),
    .A2(_01187_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06378_ (.A1(_01254_),
    .A2(_01257_),
    .B(_01258_),
    .C(_01228_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06379_ (.A1(_01229_),
    .A2(_01124_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06380_ (.A1(_01146_),
    .A2(_01260_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06381_ (.A1(_01253_),
    .A2(_01261_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06382_ (.A1(_01239_),
    .A2(_01254_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06383_ (.I(_01085_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06384_ (.I(_01088_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06385_ (.A1(_01264_),
    .A2(_01265_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06386_ (.I(_01266_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06387_ (.A1(_01213_),
    .A2(_01235_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06388_ (.A1(_01267_),
    .A2(_01254_),
    .A3(_01268_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06389_ (.A1(_01259_),
    .A2(_01262_),
    .A3(_01263_),
    .A4(_01269_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06390_ (.A1(_01251_),
    .A2(_01270_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06391_ (.A1(_01250_),
    .A2(_01271_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06392_ (.A1(_01144_),
    .A2(_01260_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06393_ (.A1(_01208_),
    .A2(_01273_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06394_ (.I(_01274_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06395_ (.A1(_01085_),
    .A2(_00701_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06396_ (.A1(_01085_),
    .A2(_00713_),
    .B(_01276_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06397_ (.A1(_01084_),
    .A2(_00881_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06398_ (.A1(_01084_),
    .A2(_00888_),
    .B(_01278_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06399_ (.I(_01279_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06400_ (.I(_00864_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06401_ (.A1(_00862_),
    .A2(_00824_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06402_ (.A1(_01084_),
    .A2(_00833_),
    .B(_01282_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06403_ (.I(_00806_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06404_ (.I(_00785_),
    .Z(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06405_ (.I(_00760_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06406_ (.I(_01006_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06407_ (.I(_00684_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06408_ (.I0(_00726_),
    .I1(_01287_),
    .S(_01288_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06409_ (.I(_00739_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06410_ (.I0(_00735_),
    .I1(_01290_),
    .S(_00684_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06411_ (.I0(_01289_),
    .I1(_01291_),
    .S(_00674_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06412_ (.A1(_01286_),
    .A2(_01292_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06413_ (.A1(_01285_),
    .A2(_01293_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06414_ (.A1(_01283_),
    .A2(_01284_),
    .A3(_01294_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06415_ (.A1(_01281_),
    .A2(_01295_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06416_ (.A1(_01280_),
    .A2(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06417_ (.A1(_01277_),
    .A2(_01297_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06418_ (.A1(_01275_),
    .A2(_01298_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06419_ (.I(_00716_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06420_ (.A1(_01236_),
    .A2(_01273_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06421_ (.I(_01283_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06422_ (.I(_01284_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06423_ (.I(_00741_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06424_ (.A1(_01303_),
    .A2(_01285_),
    .A3(_01033_),
    .A4(_01304_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06425_ (.A1(_01302_),
    .A2(_01305_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06426_ (.A1(_01281_),
    .A2(_01306_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06427_ (.A1(_01280_),
    .A2(_01307_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _06428_ (.A1(_00716_),
    .A2(_01308_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06429_ (.A1(_01300_),
    .A2(_01273_),
    .B1(_01301_),
    .B2(_01309_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06430_ (.A1(_01299_),
    .A2(_01310_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06431_ (.I(_00890_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06432_ (.A1(_01230_),
    .A2(_01125_),
    .A3(_01210_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06433_ (.I(_01313_),
    .Z(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06434_ (.I(_01314_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06435_ (.A1(_01208_),
    .A2(_01313_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06436_ (.I(_01316_),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06437_ (.A1(_00890_),
    .A2(_01307_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06438_ (.I(_01318_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06439_ (.A1(_01280_),
    .A2(_01296_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06440_ (.A1(_01275_),
    .A2(_01320_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06441_ (.A1(_01312_),
    .A2(_01315_),
    .B1(_01317_),
    .B2(_01319_),
    .C(_01321_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06442_ (.I(_01322_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06443_ (.I(_00864_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06444_ (.A1(_01324_),
    .A2(_01306_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06445_ (.A1(_01281_),
    .A2(_01295_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06446_ (.A1(_01275_),
    .A2(_01326_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06447_ (.A1(_01324_),
    .A2(_01315_),
    .B1(_01317_),
    .B2(_01325_),
    .C(_01327_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06448_ (.I(_00835_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06449_ (.I(_01329_),
    .Z(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06450_ (.A1(_01302_),
    .A2(_01305_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06451_ (.I(_01284_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06452_ (.A1(_01332_),
    .A2(_01294_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06453_ (.A1(_01329_),
    .A2(_01333_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06454_ (.A1(_01275_),
    .A2(_01334_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06455_ (.A1(_01330_),
    .A2(_01315_),
    .B1(_01317_),
    .B2(_01331_),
    .C(_01335_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06456_ (.I0(_00777_),
    .I1(_00782_),
    .S(_01288_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06457_ (.I0(_00773_),
    .I1(_01337_),
    .S(_01226_),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06458_ (.I(_01338_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06459_ (.I(_01033_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06460_ (.I(_01304_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06461_ (.A1(_01340_),
    .A2(_01341_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06462_ (.A1(_01339_),
    .A2(_01342_),
    .B(_01332_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06463_ (.A1(_01305_),
    .A2(_01343_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06464_ (.A1(_01316_),
    .A2(_01344_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06465_ (.I(_01332_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06466_ (.A1(_01136_),
    .A2(_01313_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06467_ (.A1(_01332_),
    .A2(_01294_),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06468_ (.A1(_01346_),
    .A2(_01314_),
    .B1(_01347_),
    .B2(_01348_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06469_ (.A1(_01345_),
    .A2(_01349_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06470_ (.I(_01339_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06471_ (.A1(_01285_),
    .A2(_01342_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06472_ (.A1(_01339_),
    .A2(_01293_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06473_ (.A1(_01274_),
    .A2(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06474_ (.A1(_01351_),
    .A2(_01314_),
    .B1(_01316_),
    .B2(_01352_),
    .C(_01354_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06475_ (.A1(_01293_),
    .A2(_01342_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06476_ (.A1(_01341_),
    .A2(_01313_),
    .B(_01347_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06477_ (.A1(_01356_),
    .A2(_01357_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06478_ (.I(_01292_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06479_ (.A1(_01359_),
    .A2(_01314_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06480_ (.A1(_01355_),
    .A2(_01358_),
    .A3(_01360_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06481_ (.A1(_01328_),
    .A2(_01336_),
    .A3(_01350_),
    .A4(_01361_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06482_ (.I(_01125_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06483_ (.A1(_01311_),
    .A2(_01323_),
    .A3(_01362_),
    .B1(_01255_),
    .B2(_01363_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06484_ (.A1(\as2650.debug_psl[6] ),
    .A2(_01288_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06485_ (.A1(\as2650.debug_psl[7] ),
    .A2(_01226_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06486_ (.A1(_01365_),
    .A2(_01366_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06487_ (.A1(_01230_),
    .A2(_01363_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06488_ (.A1(_01266_),
    .A2(_01367_),
    .B(_01368_),
    .C(_01220_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06489_ (.A1(_01234_),
    .A2(_01367_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06490_ (.A1(_01159_),
    .A2(_01161_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06491_ (.I(_01371_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06492_ (.A1(_01114_),
    .A2(_01125_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06493_ (.A1(_01082_),
    .A2(_01145_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06494_ (.A1(_01373_),
    .A2(_01374_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06495_ (.A1(_01264_),
    .A2(_01265_),
    .A3(_01372_),
    .A4(_01375_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06496_ (.A1(_01092_),
    .A2(_01161_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06497_ (.A1(_01264_),
    .A2(_01088_),
    .A3(_01377_),
    .A4(_01375_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06498_ (.I(_01378_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06499_ (.A1(_01221_),
    .A2(_01376_),
    .A3(_01379_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _06500_ (.A1(_01364_),
    .A2(_01369_),
    .A3(_01370_),
    .A4(_01380_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06501_ (.I(_01381_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06502_ (.I(_01382_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06503_ (.I(_01383_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06504_ (.A1(_01272_),
    .A2(_01384_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06505_ (.A1(_01207_),
    .A2(_01385_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06506_ (.I(\as2650.is_interrupt_cycle ),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06507_ (.I(_01387_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06508_ (.I(_01388_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06509_ (.I(_00983_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06510_ (.A1(_01390_),
    .A2(_01197_),
    .A3(_01200_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06511_ (.A1(_00982_),
    .A2(_01223_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06512_ (.I(_01392_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06513_ (.A1(_01171_),
    .A2(_01393_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06514_ (.I(_01394_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06515_ (.A1(_01389_),
    .A2(_01391_),
    .A3(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06516_ (.I(_01252_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06517_ (.A1(_00602_),
    .A2(_01397_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06518_ (.I(_01398_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06519_ (.I(_01399_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06520_ (.I(_01221_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06521_ (.I(_00593_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06522_ (.I(_01110_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06523_ (.A1(_00940_),
    .A2(_01219_),
    .A3(_01403_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06524_ (.I(_01371_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06525_ (.A1(_01404_),
    .A2(_01405_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06526_ (.A1(_01402_),
    .A2(_01163_),
    .A3(_01406_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06527_ (.A1(_01187_),
    .A2(_01404_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06528_ (.I(_01408_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06529_ (.A1(_01401_),
    .A2(_01407_),
    .B(_01409_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06530_ (.I(_01195_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06531_ (.A1(_01400_),
    .A2(_01410_),
    .B(_01411_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06532_ (.A1(_01079_),
    .A2(_01073_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06533_ (.A1(_01200_),
    .A2(_01412_),
    .A3(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06534_ (.A1(_01220_),
    .A2(_01404_),
    .B(_01200_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06535_ (.A1(_01402_),
    .A2(_01250_),
    .A3(_01398_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06536_ (.I(_01416_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06537_ (.A1(_01372_),
    .A2(_01415_),
    .B(_01417_),
    .C(_01186_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06538_ (.A1(_01414_),
    .A2(_01418_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06539_ (.A1(_01168_),
    .A2(_01419_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06540_ (.A1(_01249_),
    .A2(_01386_),
    .B1(_01396_),
    .B2(_01184_),
    .C(_01420_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06541_ (.I(_01209_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06542_ (.A1(_01188_),
    .A2(_01374_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06543_ (.A1(_01233_),
    .A2(_01421_),
    .A3(_01422_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06544_ (.I(_01226_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06545_ (.I(_01209_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06546_ (.I(_01373_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06547_ (.I(_01426_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06548_ (.A1(_01425_),
    .A2(_01427_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06549_ (.A1(_01424_),
    .A2(_01422_),
    .A3(_01428_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06550_ (.A1(_01390_),
    .A2(_00974_),
    .A3(_01063_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06551_ (.I(_01430_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06552_ (.A1(_01082_),
    .A2(_01103_),
    .B(_01261_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06553_ (.A1(_01083_),
    .A2(_01160_),
    .B(_01432_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06554_ (.I(_01433_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06555_ (.A1(_01190_),
    .A2(_01434_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06556_ (.A1(_01431_),
    .A2(_01435_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06557_ (.A1(_01429_),
    .A2(_01436_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06558_ (.A1(_01423_),
    .A2(_01437_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06559_ (.I(_01438_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06560_ (.I(_01439_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06561_ (.A1(_01202_),
    .A2(_01440_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06562_ (.I(_01441_),
    .Z(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06563_ (.I(_01176_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06564_ (.I(_01442_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06565_ (.I(_01443_),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06566_ (.A1(_01148_),
    .A2(_01216_),
    .A3(_01249_),
    .A4(_01385_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06567_ (.A1(_01198_),
    .A2(_01445_),
    .B(_01207_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06568_ (.I(_01196_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06569_ (.I(_01447_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06570_ (.I(\as2650.cycle[10] ),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06571_ (.A1(_01449_),
    .A2(_00977_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06572_ (.A1(_01207_),
    .A2(_01074_),
    .B(_01450_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06573_ (.I(_01255_),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06574_ (.A1(_01164_),
    .A2(_01404_),
    .A3(_01405_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06575_ (.A1(_01452_),
    .A2(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06576_ (.A1(_01400_),
    .A2(_01454_),
    .B(_01167_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06577_ (.I(_01193_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06578_ (.A1(_01221_),
    .A2(_01223_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06579_ (.A1(_01456_),
    .A2(_01457_),
    .B(_00938_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06580_ (.A1(_01423_),
    .A2(_01455_),
    .B(_01458_),
    .C(_01450_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06581_ (.A1(\as2650.cycle[11] ),
    .A2(_01074_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06582_ (.A1(_01448_),
    .A2(_01451_),
    .B(_01459_),
    .C(_01460_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06583_ (.A1(_01444_),
    .A2(_01446_),
    .A3(_01461_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06584_ (.I(_00727_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06585_ (.I(_01462_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06586_ (.I(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06587_ (.I(_01464_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06588_ (.I(_01465_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06589_ (.I(_01466_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06590_ (.I(_01467_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06591_ (.I(_01468_),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06592_ (.I(_00747_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06593_ (.I(_01469_),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06594_ (.I(_01470_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06595_ (.I(_01471_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06596_ (.I(_01472_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06597_ (.I(_01473_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06598_ (.I(_01474_),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06599_ (.I(_00770_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06600_ (.I(_01475_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06601_ (.I(_01476_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06602_ (.I(_01477_),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06603_ (.I(_01478_),
    .Z(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06604_ (.I(_01479_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06605_ (.I(_01480_),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06606_ (.I(_00793_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06607_ (.I(_01481_),
    .Z(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06608_ (.I(_01482_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06609_ (.I(_01483_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06610_ (.I(_01484_),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06611_ (.I(wb_io3_test),
    .ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06612_ (.A1(_01078_),
    .A2(_01183_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06613_ (.I(_01485_),
    .Z(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06614_ (.A1(\as2650.cycle[2] ),
    .A2(_00977_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06615_ (.I(_01486_),
    .Z(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06616_ (.I(_01172_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06617_ (.A1(\as2650.cycle[2] ),
    .A2(_01231_),
    .A3(_01216_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06618_ (.A1(_00602_),
    .A2(_01390_),
    .B(_00650_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06619_ (.A1(_01434_),
    .A2(_01490_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06620_ (.A1(_01487_),
    .A2(_01488_),
    .B1(_01489_),
    .B2(_01491_),
    .C(_01079_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06621_ (.I(_01492_),
    .ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06622_ (.I(\as2650.io_bus_we ),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06623_ (.I(\as2650.ext_io_addr[7] ),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06624_ (.I(_01494_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06625_ (.I(\as2650.ext_io_addr[6] ),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06626_ (.I(_01496_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06627_ (.A1(_01493_),
    .A2(_01495_),
    .A3(_01497_),
    .ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06628_ (.I(_01495_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06629_ (.A1(\as2650.io_bus_we ),
    .A2(_01498_),
    .A3(_01497_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06630_ (.I(_01499_),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06631_ (.A1(_01493_),
    .A2(_01498_),
    .A3(_01497_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06632_ (.A1(\as2650.io_bus_we ),
    .A2(_01495_),
    .A3(_01497_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06633_ (.I(_01500_),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06634_ (.I(_01115_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06635_ (.A1(_01486_),
    .A2(_01501_),
    .A3(_01213_),
    .A4(_01215_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06636_ (.I(_01502_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06637_ (.A1(_00989_),
    .A2(_01068_),
    .A3(_01492_),
    .A4(_01503_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06638_ (.A1(_01444_),
    .A2(_01504_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06639_ (.I(_01488_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06640_ (.A1(_01501_),
    .A2(_01216_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06641_ (.A1(_00984_),
    .A2(_01505_),
    .B1(_01506_),
    .B2(_01487_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06642_ (.A1(_01444_),
    .A2(_01491_),
    .A3(_01507_),
    .ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06643_ (.I(_01442_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06644_ (.I(_01508_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06645_ (.A1(clknet_leaf_51_wb_clk_i),
    .A2(_00989_),
    .A3(_01509_),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06646_ (.I(_01510_),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06647_ (.A1(clknet_leaf_51_wb_clk_i),
    .A2(net238),
    .A3(_01509_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06648_ (.I(_01511_),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06649_ (.A1(\web_behavior[1] ),
    .A2(clknet_leaf_141_wb_clk_i),
    .B(\web_behavior[0] ),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06650_ (.A1(\web_behavior[1] ),
    .A2(clknet_leaf_141_wb_clk_i),
    .B(\web_behavior[0] ),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06651__1 (.I(_01513_),
    .ZN(net348));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06652_ (.A1(_01512_),
    .A2(net348),
    .B(net309),
    .ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06653_ (.I(wb_debug_carry),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06654_ (.I(\as2650.debug_psl[0] ),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06655_ (.I(_01516_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06656_ (.I(_01517_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06657_ (.I(wb_debug_cc),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06658_ (.I(\as2650.debug_psl[6] ),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06659_ (.I(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06660_ (.I(\as2650.insin[6] ),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06661_ (.A1(_01522_),
    .A2(wb_debug_cc),
    .A3(_01487_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06662_ (.A1(_01519_),
    .A2(_01521_),
    .B(_01523_),
    .C(wb_debug_carry),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06663_ (.A1(_01515_),
    .A2(_01518_),
    .B(_01524_),
    .ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06664_ (.I(\as2650.debug_psl[7] ),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06665_ (.A1(\as2650.insin[6] ),
    .A2(_01519_),
    .A3(_01487_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06666_ (.A1(_01519_),
    .A2(_01525_),
    .B(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06667_ (.I(\as2650.debug_psl[5] ),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06668_ (.I(_01528_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06669_ (.I(_01529_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06670_ (.A1(_01515_),
    .A2(_01530_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06671_ (.A1(_01515_),
    .A2(_01527_),
    .B(_01531_),
    .ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06672_ (.I(_00753_),
    .ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06673_ (.I(_00800_),
    .ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06674_ (.I(_00739_),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06675_ (.I(_00756_),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06676_ (.I(_00803_),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06677_ (.I(_00849_),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06678_ (.I(_00710_),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06679_ (.A1(_01241_),
    .A2(_01149_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _06680_ (.A1(_01272_),
    .A2(_01532_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06681_ (.I(_01533_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06682_ (.A1(_01238_),
    .A2(_01256_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06683_ (.A1(_01224_),
    .A2(_01228_),
    .A3(_01267_),
    .A4(_01535_),
    .Z(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06684_ (.I(_01536_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06685_ (.A1(\as2650.chirp_ptr[1] ),
    .A2(\as2650.chirp_ptr[0] ),
    .A3(_01534_),
    .A4(_01537_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06686_ (.A1(\as2650.chirp_ptr[2] ),
    .A2(_01538_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06687_ (.I(_01539_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06688_ (.A1(_01533_),
    .A2(_01537_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06689_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01541_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06690_ (.A1(_01078_),
    .A2(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06691_ (.I(_01543_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06692_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01533_),
    .A3(_01537_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06693_ (.A1(\as2650.chirp_ptr[1] ),
    .A2(_01544_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06694_ (.A1(_01176_),
    .A2(_01545_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06695_ (.I(_01546_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06696_ (.A1(_00146_),
    .A2(_00147_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06697_ (.A1(_01542_),
    .A2(_01546_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06698_ (.A1(_01547_),
    .A2(_01548_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06699_ (.I(_01176_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06700_ (.A1(_01550_),
    .A2(_01539_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06701_ (.I(_01551_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06702_ (.I(_01552_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06703_ (.A1(_01540_),
    .A2(_00146_),
    .B1(_01549_),
    .B2(_00148_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06704_ (.A1(_01552_),
    .A2(_01547_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06705_ (.A1(_01548_),
    .A2(_01553_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06706_ (.A1(_01552_),
    .A2(_01545_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06707_ (.A1(_00148_),
    .A2(_01549_),
    .B(_01554_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06708_ (.A1(_01552_),
    .A2(_01547_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06709_ (.A1(_01551_),
    .A2(_01548_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06710_ (.A1(_00515_),
    .A2(_01555_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06711_ (.I(_01556_),
    .Z(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06712_ (.A1(_01553_),
    .A2(_01554_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06713_ (.I(_01557_),
    .Z(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06714_ (.I(_01359_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06715_ (.I(_01558_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06716_ (.I(_01503_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06717_ (.I(_01066_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06718_ (.I(_01561_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06719_ (.I(_00744_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06720_ (.I(_01563_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06721_ (.I(_01564_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06722_ (.I(_01341_),
    .Z(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06723_ (.A1(_01563_),
    .A2(_00726_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06724_ (.A1(_01565_),
    .A2(_01566_),
    .B(_01567_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06725_ (.I(_00987_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06726_ (.A1(net254),
    .A2(_01569_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06727_ (.A1(_00989_),
    .A2(_01568_),
    .B(_01570_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06728_ (.A1(_01562_),
    .A2(_01571_),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06729_ (.I(_01067_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06730_ (.I(_01503_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06731_ (.A1(net240),
    .A2(_01573_),
    .B(_01574_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06732_ (.A1(_01559_),
    .A2(_01560_),
    .B1(_01572_),
    .B2(_01575_),
    .ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06733_ (.I(_01286_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06734_ (.I(_00987_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06735_ (.I(_00747_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06736_ (.I0(_01578_),
    .I1(_00760_),
    .S(_00744_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06737_ (.I(_00987_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06738_ (.A1(net255),
    .A2(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06739_ (.A1(_01577_),
    .A2(_01579_),
    .B(_01581_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06740_ (.A1(_01562_),
    .A2(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06741_ (.A1(net247),
    .A2(_01573_),
    .B(_01574_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06742_ (.A1(_01576_),
    .A2(_01560_),
    .B1(_01583_),
    .B2(_01584_),
    .ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06743_ (.I(_01351_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06744_ (.I(_01585_),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06745_ (.I(_00770_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06746_ (.I0(_01587_),
    .I1(_01338_),
    .S(_01563_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06747_ (.I(_01588_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06748_ (.A1(net241),
    .A2(_00988_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06749_ (.A1(_01577_),
    .A2(_01589_),
    .B(_01590_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06750_ (.A1(_01562_),
    .A2(_01591_),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06751_ (.A1(net248),
    .A2(_01573_),
    .B(_01574_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06752_ (.A1(_01586_),
    .A2(_01560_),
    .B1(_01592_),
    .B2(_01593_),
    .ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06753_ (.I(_01346_),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06754_ (.I(_01594_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06755_ (.I(_01561_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06756_ (.I0(_00794_),
    .I1(_00806_),
    .S(_00744_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06757_ (.I(_01597_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06758_ (.A1(net242),
    .A2(_01569_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06759_ (.A1(_01577_),
    .A2(_01598_),
    .B(_01599_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06760_ (.A1(_01596_),
    .A2(_01600_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06761_ (.I(_01067_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06762_ (.A1(net249),
    .A2(_01602_),
    .B(_01574_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06763_ (.A1(_01595_),
    .A2(_01560_),
    .B1(_01601_),
    .B2(_01603_),
    .ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06764_ (.I(_01302_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06765_ (.I(_01604_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06766_ (.I(_01503_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06767_ (.I(_00816_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06768_ (.A1(_01564_),
    .A2(_01607_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06769_ (.A1(_01564_),
    .A2(_01329_),
    .B(_01608_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06770_ (.I(_01609_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06771_ (.A1(net243),
    .A2(_00988_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06772_ (.A1(_01577_),
    .A2(_01610_),
    .B(_01611_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06773_ (.A1(_01596_),
    .A2(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06774_ (.I(_01502_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06775_ (.A1(net250),
    .A2(_01602_),
    .B(_01614_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06776_ (.A1(_01605_),
    .A2(_01606_),
    .B1(_01613_),
    .B2(_01615_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06777_ (.A1(_00851_),
    .A2(_00863_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06778_ (.I(_01616_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06779_ (.I(_01617_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06780_ (.A1(_01564_),
    .A2(_00855_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06781_ (.A1(_01565_),
    .A2(_01281_),
    .B(_01619_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06782_ (.A1(net244),
    .A2(_01569_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06783_ (.A1(_01580_),
    .A2(_01620_),
    .B(_01621_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06784_ (.A1(_01596_),
    .A2(_01622_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06785_ (.A1(net251),
    .A2(_01602_),
    .B(_01614_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06786_ (.A1(_01618_),
    .A2(_01606_),
    .B1(_01623_),
    .B2(_01624_),
    .ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06787_ (.I(_01280_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06788_ (.I(_01625_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06789_ (.I(_01626_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06790_ (.I(_01028_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06791_ (.I(_01628_),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06792_ (.A1(_01628_),
    .A2(_01279_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06793_ (.A1(_01629_),
    .A2(_01013_),
    .B(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06794_ (.I(_01631_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06795_ (.A1(net245),
    .A2(_00988_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06796_ (.A1(_01580_),
    .A2(_01632_),
    .B(_01633_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06797_ (.A1(_01596_),
    .A2(_01634_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06798_ (.A1(net252),
    .A2(_01602_),
    .B(_01614_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06799_ (.A1(_01627_),
    .A2(_01606_),
    .B1(_01635_),
    .B2(_01636_),
    .ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06800_ (.I(_01277_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06801_ (.I(_01637_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06802_ (.I(_00693_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06803_ (.A1(_01565_),
    .A2(_01639_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06804_ (.A1(_01565_),
    .A2(_00716_),
    .B(_01640_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06805_ (.I(_01641_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06806_ (.A1(net246),
    .A2(_01569_),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06807_ (.A1(_01580_),
    .A2(_01642_),
    .B(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06808_ (.A1(_01561_),
    .A2(_01644_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06809_ (.A1(net253),
    .A2(_01068_),
    .B(_01614_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06810_ (.A1(_01638_),
    .A2(_01606_),
    .B1(_01645_),
    .B2(_01646_),
    .ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06811_ (.I(_01177_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06812_ (.I(_01647_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06813_ (.A1(_00983_),
    .A2(_01179_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06814_ (.I(_01649_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06815_ (.I(_01650_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06816_ (.A1(_01648_),
    .A2(_00601_),
    .A3(_01651_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06817_ (.I(_01431_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06818_ (.I(_01653_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06819_ (.I(_01654_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06820_ (.A1(_01220_),
    .A2(_01406_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06821_ (.I(_01656_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06822_ (.A1(_01417_),
    .A2(_01655_),
    .A3(_01657_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06823_ (.I(_01077_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06824_ (.I(_01659_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06825_ (.I(_01660_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06826_ (.I(_01661_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06827_ (.A1(_01652_),
    .A2(_01658_),
    .B(_01662_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06828_ (.I(net105),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06829_ (.A1(net104),
    .A2(net71),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06830_ (.A1(wb_feedback_delay),
    .A2(_01664_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06831_ (.I(_01665_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06832_ (.I(net70),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06833_ (.A1(net427),
    .A2(_01667_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06834_ (.I(net67),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06835_ (.I(_01669_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06836_ (.A1(_01670_),
    .A2(net68),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06837_ (.A1(net66),
    .A2(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06838_ (.A1(_01663_),
    .A2(_01666_),
    .A3(_01668_),
    .A4(_01672_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06839_ (.I(_01673_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06840_ (.I(_01674_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06841_ (.I0(net72),
    .I1(net122),
    .S(_01675_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06842_ (.I(_01676_),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06843_ (.I0(net83),
    .I1(net129),
    .S(_01675_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06844_ (.I(_01677_),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06845_ (.I0(net94),
    .I1(net130),
    .S(_01675_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06846_ (.I(_01678_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06847_ (.I0(net97),
    .I1(net131),
    .S(_01675_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06848_ (.I(_01679_),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06849_ (.I(_01674_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06850_ (.I0(net98),
    .I1(net132),
    .S(_01680_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06851_ (.I(_01681_),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06852_ (.I0(net99),
    .I1(net133),
    .S(_01680_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06853_ (.I(_01682_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06854_ (.I0(net100),
    .I1(net134),
    .S(_01680_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06855_ (.I(_01683_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06856_ (.I0(net101),
    .I1(net135),
    .S(_01680_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06857_ (.I(_01684_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06858_ (.I(_01674_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06859_ (.I0(net102),
    .I1(net136),
    .S(_01685_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06860_ (.I(_01686_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06861_ (.I0(net103),
    .I1(net137),
    .S(_01685_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06862_ (.I(_01687_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06863_ (.I0(net73),
    .I1(net123),
    .S(_01685_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06864_ (.I(_01688_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06865_ (.I0(net74),
    .I1(net124),
    .S(_01685_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06866_ (.I(_01689_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06867_ (.I(_01674_),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06868_ (.I0(net75),
    .I1(net125),
    .S(_01690_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06869_ (.I(_01691_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06870_ (.I0(net76),
    .I1(net126),
    .S(_01690_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06871_ (.I(_01692_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06872_ (.I0(net77),
    .I1(net127),
    .S(_01690_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06873_ (.I(_01693_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06874_ (.I0(net78),
    .I1(net128),
    .S(_01690_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06875_ (.I(_01694_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06876_ (.I(_01673_),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06877_ (.I(_01695_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06878_ (.I0(net79),
    .I1(net106),
    .S(_01696_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06879_ (.I(_01697_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06880_ (.I0(net80),
    .I1(net113),
    .S(_01696_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06881_ (.I(_01698_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06882_ (.I0(net81),
    .I1(net114),
    .S(_01696_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06883_ (.I(_01699_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06884_ (.I0(net82),
    .I1(net115),
    .S(_01696_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06885_ (.I(_01700_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06886_ (.I(_01695_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06887_ (.I0(net84),
    .I1(net116),
    .S(_01701_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06888_ (.I(_01702_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06889_ (.I0(net85),
    .I1(net117),
    .S(_01701_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06890_ (.I(_01703_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06891_ (.I0(net86),
    .I1(net118),
    .S(_01701_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06892_ (.I(_01704_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06893_ (.I0(net87),
    .I1(net119),
    .S(_01701_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06894_ (.I(_01705_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06895_ (.I(_01695_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06896_ (.I0(net88),
    .I1(net120),
    .S(_01706_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06897_ (.I(_01707_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06898_ (.I0(net89),
    .I1(net121),
    .S(_01706_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06899_ (.I(_01708_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06900_ (.I0(net90),
    .I1(net107),
    .S(_01706_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06901_ (.I(_01709_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06902_ (.I0(net91),
    .I1(net108),
    .S(_01706_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06903_ (.I(_01710_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06904_ (.I(_01695_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06905_ (.I0(net92),
    .I1(net109),
    .S(_01711_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06906_ (.I(_01712_),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06907_ (.I0(net93),
    .I1(net110),
    .S(_01711_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06908_ (.I(_01713_),
    .Z(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06909_ (.I0(net95),
    .I1(net111),
    .S(_01711_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06910_ (.I(_01714_),
    .Z(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06911_ (.I0(net96),
    .I1(net112),
    .S(_01711_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06912_ (.I(_01715_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06913_ (.I(net69),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06914_ (.I(_01667_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06915_ (.A1(_01663_),
    .A2(_01716_),
    .A3(_01717_),
    .A4(_01666_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06916_ (.I(_01718_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06917_ (.I(_01719_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06918_ (.A1(net102),
    .A2(_01719_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06919_ (.I(net66),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06920_ (.I(_01722_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06921_ (.I(_01723_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06922_ (.A1(_00663_),
    .A2(_01720_),
    .B(_01721_),
    .C(_01724_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06923_ (.I(_01722_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06924_ (.I(net68),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06925_ (.A1(_01669_),
    .A2(_01726_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06926_ (.I(_01727_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06927_ (.A1(_01663_),
    .A2(_01666_),
    .A3(_01668_),
    .A4(_01728_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06928_ (.A1(_01725_),
    .A2(_01729_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06929_ (.I0(net159),
    .I1(net72),
    .S(_01730_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06930_ (.I(_01731_),
    .Z(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06931_ (.I0(net160),
    .I1(net83),
    .S(_01730_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06932_ (.I(_01732_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06933_ (.I0(net161),
    .I1(net94),
    .S(_01730_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06934_ (.I(_01733_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06935_ (.I(_01722_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06936_ (.I(_01734_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06937_ (.I(_01735_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06938_ (.A1(_01736_),
    .A2(wb_feedback_delay),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06939_ (.I(_01737_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06940_ (.A1(wb_feedback_delay),
    .A2(_01664_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06941_ (.I(_01738_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06942_ (.I(_01739_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06943_ (.A1(net266),
    .A2(_01740_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06944_ (.I(net70),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06945_ (.I(_01742_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06946_ (.I(_01743_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06947_ (.I(net69),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06948_ (.I(_01745_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06949_ (.A1(_01726_),
    .A2(_01746_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06950_ (.A1(_01670_),
    .A2(net122),
    .B1(net159),
    .B2(_01728_),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06951_ (.A1(_01746_),
    .A2(_01518_),
    .B1(_01747_),
    .B2(_01748_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06952_ (.I(_01743_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06953_ (.I(\wb_counter[0] ),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06954_ (.A1(_01750_),
    .A2(_01751_),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06955_ (.I(_01665_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06956_ (.A1(_01744_),
    .A2(_01749_),
    .B(_01752_),
    .C(_01753_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06957_ (.I(_01722_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06958_ (.I(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06959_ (.A1(_01741_),
    .A2(_01754_),
    .B(_01756_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06960_ (.A1(net277),
    .A2(_01740_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06961_ (.I(\as2650.debug_psl[1] ),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06962_ (.I(_01758_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06963_ (.I(_01759_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06964_ (.A1(net67),
    .A2(net160),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06965_ (.I(_01716_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06966_ (.A1(_01670_),
    .A2(net129),
    .B(_01762_),
    .C(_01726_),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06967_ (.A1(_01746_),
    .A2(_01760_),
    .B1(_01761_),
    .B2(_01763_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06968_ (.I(\wb_counter[1] ),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06969_ (.A1(_01750_),
    .A2(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06970_ (.A1(_01744_),
    .A2(net476),
    .B(_01766_),
    .C(_01753_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06971_ (.A1(_01757_),
    .A2(_01767_),
    .B(_01756_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06972_ (.A1(net288),
    .A2(_01740_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06973_ (.I(\as2650.debug_psl[2] ),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06974_ (.I(_01769_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06975_ (.A1(net67),
    .A2(net161),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06976_ (.A1(_01670_),
    .A2(net130),
    .B(_01762_),
    .C(_01726_),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06977_ (.A1(_01746_),
    .A2(_01770_),
    .B1(_01771_),
    .B2(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06978_ (.I(_01667_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06979_ (.I(_01774_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06980_ (.I(\wb_counter[2] ),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06981_ (.A1(_01775_),
    .A2(_01776_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06982_ (.A1(_01744_),
    .A2(_01773_),
    .B(_01777_),
    .C(_01753_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06983_ (.A1(_01768_),
    .A2(_01778_),
    .B(_01756_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06984_ (.I(_01723_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06985_ (.I(_01738_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06986_ (.I(_01780_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06987_ (.I(\wb_counter[3] ),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06988_ (.I(_01671_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06989_ (.I(_01783_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06990_ (.A1(net69),
    .A2(_01727_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06991_ (.I(_01785_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06992_ (.I(_01786_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06993_ (.A1(net131),
    .A2(_01784_),
    .B(_01787_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06994_ (.I(_01745_),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06995_ (.I(\as2650.debug_psl[3] ),
    .Z(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06996_ (.I(_01790_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06997_ (.I(_01791_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06998_ (.I(_01742_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06999_ (.A1(_01789_),
    .A2(_01792_),
    .B(_01793_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07000_ (.I(_01738_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07001_ (.A1(_01775_),
    .A2(_01782_),
    .B1(_01788_),
    .B2(_01794_),
    .C(_01795_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07002_ (.A1(net291),
    .A2(_01781_),
    .B(_01796_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07003_ (.A1(_01779_),
    .A2(_01797_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07004_ (.I(_01780_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07005_ (.I(\wb_counter[4] ),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07006_ (.I(_01783_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07007_ (.A1(net132),
    .A2(_01800_),
    .B(_01787_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07008_ (.I(_00707_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07009_ (.I(_01802_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07010_ (.I(_01803_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07011_ (.I(_01716_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07012_ (.I(_01774_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07013_ (.A1(_01804_),
    .A2(_01805_),
    .B(_01806_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07014_ (.A1(_01775_),
    .A2(_01799_),
    .B1(_01801_),
    .B2(_01807_),
    .C(_01795_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07015_ (.A1(net292),
    .A2(_01798_),
    .B(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07016_ (.A1(_01779_),
    .A2(_01809_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07017_ (.I(_01755_),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07018_ (.I(\wb_counter[5] ),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07019_ (.A1(net133),
    .A2(_01800_),
    .B(_01787_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07020_ (.A1(_01789_),
    .A2(_01530_),
    .B(_01806_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07021_ (.I(_01738_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07022_ (.I(_01814_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07023_ (.A1(_01775_),
    .A2(_01811_),
    .B1(_01812_),
    .B2(_01813_),
    .C(_01815_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07024_ (.A1(net293),
    .A2(_01798_),
    .B(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07025_ (.A1(_01810_),
    .A2(_01817_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07026_ (.I(_01743_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07027_ (.I(\wb_counter[6] ),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07028_ (.A1(net134),
    .A2(_01800_),
    .B(_01787_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07029_ (.A1(_01789_),
    .A2(_01521_),
    .B(_01806_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07030_ (.A1(_01818_),
    .A2(_01819_),
    .B1(_01820_),
    .B2(_01821_),
    .C(_01815_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07031_ (.A1(net294),
    .A2(_01798_),
    .B(_01822_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07032_ (.A1(_01810_),
    .A2(_01823_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07033_ (.I(\wb_counter[7] ),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07034_ (.I(_01786_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07035_ (.A1(net135),
    .A2(_01800_),
    .B(_01825_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07036_ (.A1(_01789_),
    .A2(_01525_),
    .B(_01806_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07037_ (.A1(_01818_),
    .A2(_01824_),
    .B1(_01826_),
    .B2(_01827_),
    .C(_01815_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07038_ (.A1(net295),
    .A2(_01798_),
    .B(_01828_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07039_ (.A1(_01810_),
    .A2(_01829_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07040_ (.I(_01780_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07041_ (.I(\wb_counter[8] ),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07042_ (.I(_01783_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07043_ (.A1(net136),
    .A2(_01832_),
    .B(_01825_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07044_ (.I(_01745_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07045_ (.I(\as2650.debug_psu[0] ),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07046_ (.I(_01835_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07047_ (.I(_01836_),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07048_ (.I(_01837_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07049_ (.I(_01838_),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07050_ (.I(_01839_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07051_ (.I(_01840_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07052_ (.I(_01841_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07053_ (.I(_01842_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07054_ (.I(_01843_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07055_ (.I(_01774_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07056_ (.A1(_01834_),
    .A2(_01844_),
    .B(_01845_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07057_ (.A1(_01818_),
    .A2(_01831_),
    .B1(_01833_),
    .B2(_01846_),
    .C(_01815_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07058_ (.A1(net296),
    .A2(_01830_),
    .B(_01847_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07059_ (.A1(_01810_),
    .A2(_01848_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07060_ (.I(_01755_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07061_ (.I(\wb_counter[9] ),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07062_ (.A1(net137),
    .A2(_01832_),
    .B(_01825_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07063_ (.I(\as2650.debug_psu[1] ),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07064_ (.I(_01852_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07065_ (.A1(_01834_),
    .A2(_01853_),
    .B(_01845_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07066_ (.I(_01814_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07067_ (.A1(_01818_),
    .A2(_01850_),
    .B1(_01851_),
    .B2(_01854_),
    .C(_01855_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07068_ (.A1(net297),
    .A2(_01830_),
    .B(_01856_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07069_ (.A1(_01849_),
    .A2(_01857_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07070_ (.I(_01743_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07071_ (.I(\wb_counter[10] ),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07072_ (.A1(net123),
    .A2(_01832_),
    .B(_01825_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07073_ (.I(\as2650.debug_psu[2] ),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07074_ (.I(_01861_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07075_ (.I(_01862_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07076_ (.A1(_01834_),
    .A2(_01863_),
    .B(_01845_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07077_ (.A1(_01858_),
    .A2(_01859_),
    .B1(_01860_),
    .B2(_01864_),
    .C(_01855_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07078_ (.A1(net267),
    .A2(_01830_),
    .B(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07079_ (.A1(_01849_),
    .A2(_01866_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07080_ (.I(\wb_counter[11] ),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07081_ (.I(_01785_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07082_ (.A1(net124),
    .A2(_01832_),
    .B(_01868_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07083_ (.I(\as2650.debug_psu[3] ),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07084_ (.I(_01870_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07085_ (.A1(_01834_),
    .A2(_01871_),
    .B(_01845_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07086_ (.A1(_01858_),
    .A2(_01867_),
    .B1(_01869_),
    .B2(_01872_),
    .C(_01855_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07087_ (.A1(net268),
    .A2(_01830_),
    .B(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07088_ (.A1(_01849_),
    .A2(_01874_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07089_ (.I(_01780_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07090_ (.I(\wb_counter[12] ),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07091_ (.I(_01783_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07092_ (.A1(net125),
    .A2(_01877_),
    .B(_01868_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07093_ (.I(\as2650.debug_psu[4] ),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07094_ (.I(_01774_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07095_ (.A1(_01805_),
    .A2(_01879_),
    .B(_01880_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07096_ (.A1(_01858_),
    .A2(_01876_),
    .B1(_01878_),
    .B2(_01881_),
    .C(_01855_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07097_ (.A1(net269),
    .A2(_01875_),
    .B(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07098_ (.A1(_01849_),
    .A2(_01883_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07099_ (.I(_01755_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07100_ (.I(\wb_counter[13] ),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07101_ (.A1(net126),
    .A2(_01877_),
    .B(_01868_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07102_ (.I(\as2650.debug_psu[5] ),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07103_ (.A1(_01887_),
    .A2(_01762_),
    .B(_01880_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07104_ (.I(_01814_),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07105_ (.A1(_01858_),
    .A2(_01885_),
    .B1(_01886_),
    .B2(_01888_),
    .C(_01889_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07106_ (.A1(net270),
    .A2(_01875_),
    .B(_01890_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07107_ (.A1(_01884_),
    .A2(_01891_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07108_ (.I(\wb_counter[14] ),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07109_ (.A1(net127),
    .A2(_01877_),
    .B(_01868_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07110_ (.I(net181),
    .Z(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07111_ (.A1(_01805_),
    .A2(_01894_),
    .B(_01880_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07112_ (.A1(_01793_),
    .A2(_01892_),
    .B1(_01893_),
    .B2(_01895_),
    .C(_01889_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07113_ (.A1(net271),
    .A2(_01875_),
    .B(_01896_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07114_ (.A1(_01884_),
    .A2(_01897_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07115_ (.I(\wb_counter[15] ),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07116_ (.A1(net128),
    .A2(_01877_),
    .B(_01786_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07117_ (.I(\as2650.debug_psu[7] ),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07118_ (.A1(_01805_),
    .A2(_01900_),
    .B(_01880_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07119_ (.A1(_01793_),
    .A2(_01898_),
    .B1(_01899_),
    .B2(_01901_),
    .C(_01889_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07120_ (.A1(net272),
    .A2(_01875_),
    .B(_01902_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07121_ (.A1(_01884_),
    .A2(_01903_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07122_ (.I(\wb_counter[16] ),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07123_ (.I(_01671_),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07124_ (.A1(net106),
    .A2(_01905_),
    .B(_01786_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07125_ (.I(_01742_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07126_ (.A1(net239),
    .A2(_01762_),
    .B(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07127_ (.A1(_01793_),
    .A2(_01904_),
    .B1(_01906_),
    .B2(_01908_),
    .C(_01889_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07128_ (.A1(net273),
    .A2(_01740_),
    .B(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07129_ (.A1(_01884_),
    .A2(_01910_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07130_ (.I(net274),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07131_ (.I(_01814_),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07132_ (.I(_01912_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07133_ (.I(_01905_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07134_ (.A1(_01716_),
    .A2(_01742_),
    .A3(_01728_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07135_ (.I(_01915_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07136_ (.A1(net113),
    .A2(_01914_),
    .B(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07137_ (.I(_01739_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07138_ (.A1(_01744_),
    .A2(\wb_counter[17] ),
    .B(_01918_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07139_ (.I(_01723_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07140_ (.A1(_01911_),
    .A2(_01913_),
    .B1(_01917_),
    .B2(_01919_),
    .C(_01920_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07141_ (.I(net275),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07142_ (.A1(net114),
    .A2(_01914_),
    .B(_01916_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07143_ (.I(_01907_),
    .Z(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07144_ (.A1(_01923_),
    .A2(\wb_counter[18] ),
    .B(_01918_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07145_ (.A1(_01921_),
    .A2(_01913_),
    .B1(_01922_),
    .B2(_01924_),
    .C(_01920_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07146_ (.I(net276),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07147_ (.I(_01668_),
    .Z(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07148_ (.A1(net115),
    .A2(_01914_),
    .B(_01926_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07149_ (.A1(_01923_),
    .A2(\wb_counter[19] ),
    .B(_01918_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07150_ (.A1(_01925_),
    .A2(_01913_),
    .B1(_01927_),
    .B2(_01928_),
    .C(_01920_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07151_ (.I(net278),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07152_ (.A1(net116),
    .A2(_01914_),
    .B(_01916_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07153_ (.A1(_01923_),
    .A2(\wb_counter[20] ),
    .B(_01918_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07154_ (.I(_01725_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07155_ (.A1(_01929_),
    .A2(_01913_),
    .B1(_01930_),
    .B2(_01931_),
    .C(_01932_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07156_ (.I(net279),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07157_ (.I(_01795_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07158_ (.I(_01905_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07159_ (.A1(net117),
    .A2(_01935_),
    .B(_01916_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07160_ (.I(_01739_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07161_ (.A1(_01923_),
    .A2(\wb_counter[21] ),
    .B(_01937_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07162_ (.A1(_01933_),
    .A2(_01934_),
    .B1(_01936_),
    .B2(_01938_),
    .C(_01932_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07163_ (.I(net280),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07164_ (.I(_01915_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07165_ (.A1(net118),
    .A2(_01935_),
    .B(_01940_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07166_ (.I(_01907_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07167_ (.A1(_01942_),
    .A2(\wb_counter[22] ),
    .B(_01937_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07168_ (.A1(_01939_),
    .A2(_01934_),
    .B1(_01941_),
    .B2(_01943_),
    .C(_01932_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07169_ (.I(net281),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07170_ (.A1(net119),
    .A2(_01935_),
    .B(_01940_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07171_ (.A1(_01942_),
    .A2(\wb_counter[23] ),
    .B(_01937_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07172_ (.A1(_01944_),
    .A2(_01934_),
    .B1(_01945_),
    .B2(_01946_),
    .C(_01932_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07173_ (.I(net282),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07174_ (.A1(net120),
    .A2(_01935_),
    .B(_01926_),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07175_ (.A1(_01942_),
    .A2(\wb_counter[24] ),
    .B(_01937_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07176_ (.I(_01725_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07177_ (.A1(_01947_),
    .A2(_01934_),
    .B1(_01948_),
    .B2(_01949_),
    .C(_01950_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07178_ (.I(net283),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07179_ (.I(_01795_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07180_ (.I(_01905_),
    .Z(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07181_ (.A1(net121),
    .A2(_01953_),
    .B(_01940_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07182_ (.I(_01739_),
    .Z(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07183_ (.A1(_01942_),
    .A2(\wb_counter[25] ),
    .B(_01955_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07184_ (.A1(_01951_),
    .A2(_01952_),
    .B1(_01954_),
    .B2(_01956_),
    .C(_01950_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07185_ (.I(net284),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07186_ (.A1(net107),
    .A2(_01953_),
    .B(_01940_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07187_ (.I(_01907_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07188_ (.A1(_01959_),
    .A2(\wb_counter[26] ),
    .B(_01955_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07189_ (.A1(_01957_),
    .A2(_01952_),
    .B1(_01958_),
    .B2(_01960_),
    .C(_01950_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07190_ (.I(net285),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07191_ (.A1(net108),
    .A2(_01953_),
    .B(_01915_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07192_ (.A1(_01959_),
    .A2(\wb_counter[27] ),
    .B(_01955_),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07193_ (.A1(_01961_),
    .A2(_01952_),
    .B1(_01962_),
    .B2(_01963_),
    .C(_01950_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07194_ (.I(net286),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07195_ (.A1(net109),
    .A2(_01953_),
    .B(_01926_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07196_ (.A1(_01959_),
    .A2(\wb_counter[28] ),
    .B(_01955_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07197_ (.I(_01725_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07198_ (.A1(_01964_),
    .A2(_01952_),
    .B1(_01965_),
    .B2(_01966_),
    .C(_01967_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07199_ (.I(net287),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07200_ (.A1(net110),
    .A2(_01784_),
    .B(_01926_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07201_ (.A1(_01959_),
    .A2(\wb_counter[29] ),
    .B(_01912_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07202_ (.A1(_01968_),
    .A2(_01781_),
    .B1(_01969_),
    .B2(_01970_),
    .C(_01967_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07203_ (.I(net289),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07204_ (.A1(net111),
    .A2(_01784_),
    .B(_01915_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07205_ (.A1(_01750_),
    .A2(\wb_counter[30] ),
    .B(_01912_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07206_ (.A1(_01971_),
    .A2(_01781_),
    .B1(_01972_),
    .B2(_01973_),
    .C(_01967_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07207_ (.I(net290),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _07208_ (.I(\as2650.wb_hidden_rom_enable ),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07209_ (.A1(_01975_),
    .A2(_01728_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07210_ (.A1(net112),
    .A2(_01784_),
    .B(_01976_),
    .C(_01668_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07211_ (.A1(_01750_),
    .A2(\wb_counter[31] ),
    .B(_01912_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07212_ (.A1(_01974_),
    .A2(_01781_),
    .B1(_01977_),
    .B2(_01978_),
    .C(_01967_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07213_ (.A1(_01724_),
    .A2(net441),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07214_ (.A1(_01519_),
    .A2(_01720_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _07215_ (.A1(_01663_),
    .A2(_01745_),
    .A3(_01717_),
    .A4(_01753_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07216_ (.I(_01980_),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07217_ (.A1(net72),
    .A2(_01981_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07218_ (.A1(_01979_),
    .A2(net365),
    .B(_01756_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07219_ (.A1(_01515_),
    .A2(_01720_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07220_ (.A1(net83),
    .A2(_01981_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07221_ (.I(_01723_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07222_ (.A1(_01983_),
    .A2(net362),
    .B(_01985_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07223_ (.I(_01718_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07224_ (.A1(\web_behavior[0] ),
    .A2(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07225_ (.A1(net94),
    .A2(_01981_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07226_ (.A1(_01987_),
    .A2(net359),
    .B(_01985_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07227_ (.A1(\web_behavior[1] ),
    .A2(_01986_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07228_ (.A1(net97),
    .A2(_01981_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07229_ (.A1(_01989_),
    .A2(net356),
    .B(_01985_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07230_ (.A1(wb_reset_override_en),
    .A2(_01986_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07231_ (.A1(net98),
    .A2(_01980_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07232_ (.A1(_01991_),
    .A2(net372),
    .B(_01985_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07233_ (.A1(wb_reset_override),
    .A2(_01986_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07234_ (.A1(net99),
    .A2(_01980_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07235_ (.A1(_01993_),
    .A2(net420),
    .B(_01779_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07236_ (.A1(net100),
    .A2(_01719_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07237_ (.A1(net165),
    .A2(_01720_),
    .B(_01995_),
    .C(_01724_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07238_ (.A1(net182),
    .A2(_01719_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07239_ (.A1(net101),
    .A2(_01980_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07240_ (.A1(_01996_),
    .A2(net395),
    .B(_01779_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07241_ (.A1(net96),
    .A2(_01729_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07242_ (.A1(_01975_),
    .A2(net437),
    .B(_01998_),
    .C(_01724_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07243_ (.A1(net105),
    .A2(_01667_),
    .A3(_01666_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07244_ (.I(_01999_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07245_ (.I(_02000_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07246_ (.I(_01999_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07247_ (.I(_02002_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07248_ (.A1(net72),
    .A2(_02003_),
    .B(_01736_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07249_ (.A1(\wb_counter[0] ),
    .A2(_02001_),
    .B(_02004_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07250_ (.A1(_01751_),
    .A2(\wb_counter[1] ),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07251_ (.A1(net83),
    .A2(_02003_),
    .B(_01736_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07252_ (.A1(_02001_),
    .A2(_02005_),
    .B(_02006_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07253_ (.A1(\wb_counter[0] ),
    .A2(\wb_counter[1] ),
    .A3(\wb_counter[2] ),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07254_ (.A1(_01751_),
    .A2(_01765_),
    .B(_01776_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07255_ (.A1(_02007_),
    .A2(_02008_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07256_ (.A1(net94),
    .A2(_02003_),
    .B(_01736_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07257_ (.A1(_02001_),
    .A2(_02009_),
    .B(_02010_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07258_ (.I(_02000_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07259_ (.A1(\wb_counter[3] ),
    .A2(_02007_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07260_ (.A1(net97),
    .A2(_02000_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07261_ (.A1(_02011_),
    .A2(_02012_),
    .B(_02013_),
    .C(_01920_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07262_ (.A1(_01782_),
    .A2(_02007_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07263_ (.A1(_01799_),
    .A2(_02014_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07264_ (.I(_01735_),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07265_ (.A1(net98),
    .A2(_02003_),
    .B(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07266_ (.A1(_02001_),
    .A2(_02015_),
    .B(_02017_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07267_ (.I(_01999_),
    .Z(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07268_ (.I(_02018_),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07269_ (.I(_02019_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07270_ (.A1(\wb_counter[4] ),
    .A2(_02014_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07271_ (.A1(_01811_),
    .A2(_02021_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07272_ (.A1(\wb_counter[4] ),
    .A2(\wb_counter[5] ),
    .A3(_02014_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07273_ (.A1(_02022_),
    .A2(_02023_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07274_ (.I(_02002_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07275_ (.A1(net99),
    .A2(_02025_),
    .B(_02016_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07276_ (.A1(_02020_),
    .A2(_02024_),
    .B(_02026_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07277_ (.A1(_01819_),
    .A2(_02023_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07278_ (.A1(_01819_),
    .A2(_02023_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07279_ (.A1(_02027_),
    .A2(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07280_ (.A1(net100),
    .A2(_02025_),
    .B(_02016_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07281_ (.A1(_02020_),
    .A2(_02029_),
    .B(_02030_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07282_ (.A1(\wb_counter[7] ),
    .A2(_02028_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07283_ (.A1(net101),
    .A2(_02025_),
    .B(_02016_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07284_ (.A1(_02020_),
    .A2(_02031_),
    .B(_02032_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07285_ (.A1(_01824_),
    .A2(_02028_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07286_ (.A1(_01831_),
    .A2(_02033_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07287_ (.I(_01735_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07288_ (.A1(net102),
    .A2(_02025_),
    .B(_02035_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07289_ (.A1(_02020_),
    .A2(_02034_),
    .B(_02036_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07290_ (.I(_01999_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07291_ (.I(_02037_),
    .Z(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07292_ (.A1(_01824_),
    .A2(_01831_),
    .A3(_02028_),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07293_ (.A1(_01850_),
    .A2(_02039_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07294_ (.I(_02002_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07295_ (.A1(net103),
    .A2(_02041_),
    .B(_02035_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07296_ (.A1(_02038_),
    .A2(_02040_),
    .B(_02042_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07297_ (.A1(\wb_counter[9] ),
    .A2(_02039_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07298_ (.A1(\wb_counter[10] ),
    .A2(_02043_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07299_ (.A1(net73),
    .A2(_02041_),
    .B(_02035_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07300_ (.A1(_02038_),
    .A2(_02044_),
    .B(net414),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07301_ (.A1(_01859_),
    .A2(_02043_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07302_ (.A1(_01867_),
    .A2(_02046_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07303_ (.A1(net74),
    .A2(_02041_),
    .B(_02035_),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07304_ (.A1(_02038_),
    .A2(_02047_),
    .B(net417),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07305_ (.A1(\wb_counter[11] ),
    .A2(\wb_counter[12] ),
    .A3(_02046_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07306_ (.A1(\wb_counter[11] ),
    .A2(_02046_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07307_ (.A1(_01876_),
    .A2(_02050_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07308_ (.A1(_02049_),
    .A2(_02051_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07309_ (.I(_01735_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07310_ (.A1(net75),
    .A2(_02041_),
    .B(_02053_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07311_ (.A1(_02038_),
    .A2(_02052_),
    .B(net402),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07312_ (.I(_02037_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07313_ (.A1(\wb_counter[13] ),
    .A2(_02049_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07314_ (.I(_02002_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07315_ (.A1(net76),
    .A2(_02057_),
    .B(_02053_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07316_ (.A1(_02055_),
    .A2(_02056_),
    .B(net408),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07317_ (.A1(_01885_),
    .A2(_02049_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07318_ (.A1(_01892_),
    .A2(_02059_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07319_ (.A1(net398),
    .A2(_02057_),
    .B(_02053_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07320_ (.A1(_02055_),
    .A2(_02060_),
    .B(net399),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07321_ (.A1(\wb_counter[14] ),
    .A2(\wb_counter[15] ),
    .A3(_02059_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07322_ (.A1(\wb_counter[14] ),
    .A2(_02059_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07323_ (.A1(_01898_),
    .A2(_02063_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07324_ (.A1(_02062_),
    .A2(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07325_ (.A1(net383),
    .A2(_02057_),
    .B(_02053_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07326_ (.A1(_02055_),
    .A2(_02065_),
    .B(net384),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07327_ (.A1(\wb_counter[16] ),
    .A2(_02062_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07328_ (.I(_01734_),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07329_ (.I(_02068_),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07330_ (.A1(net379),
    .A2(_02057_),
    .B(_02069_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07331_ (.A1(_02055_),
    .A2(_02067_),
    .B(net380),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07332_ (.I(_02037_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07333_ (.A1(_01904_),
    .A2(_02062_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07334_ (.A1(\wb_counter[17] ),
    .A2(_02072_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07335_ (.I(_02018_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07336_ (.A1(net391),
    .A2(_02074_),
    .B(_02069_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07337_ (.A1(_02071_),
    .A2(_02073_),
    .B(net392),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07338_ (.A1(\wb_counter[17] ),
    .A2(_02072_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07339_ (.A1(\wb_counter[18] ),
    .A2(_02076_),
    .Z(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07340_ (.A1(net387),
    .A2(_02074_),
    .B(_02069_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07341_ (.A1(_02071_),
    .A2(_02077_),
    .B(net388),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07342_ (.A1(\wb_counter[17] ),
    .A2(\wb_counter[18] ),
    .A3(_02072_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07343_ (.A1(\wb_counter[19] ),
    .A2(_02079_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07344_ (.A1(net368),
    .A2(_02074_),
    .B(_02069_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07345_ (.A1(_02071_),
    .A2(_02080_),
    .B(net369),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07346_ (.I(\wb_counter[19] ),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07347_ (.A1(_02082_),
    .A2(_02079_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07348_ (.A1(\wb_counter[20] ),
    .A2(_02083_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07349_ (.I(_02068_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07350_ (.A1(net375),
    .A2(_02074_),
    .B(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07351_ (.A1(_02071_),
    .A2(_02084_),
    .B(net376),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07352_ (.I(_02037_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07353_ (.A1(\wb_counter[20] ),
    .A2(_02083_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07354_ (.A1(\wb_counter[21] ),
    .A2(_02088_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07355_ (.I(_02018_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07356_ (.A1(net85),
    .A2(_02090_),
    .B(_02085_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07357_ (.A1(_02087_),
    .A2(_02089_),
    .B(_02091_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07358_ (.A1(\wb_counter[20] ),
    .A2(\wb_counter[21] ),
    .A3(_02083_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07359_ (.A1(\wb_counter[22] ),
    .A2(_02092_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07360_ (.A1(net86),
    .A2(_02090_),
    .B(_02085_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07361_ (.A1(_02087_),
    .A2(_02093_),
    .B(_02094_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07362_ (.I(\wb_counter[22] ),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07363_ (.A1(_02095_),
    .A2(_02092_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07364_ (.A1(\wb_counter[23] ),
    .A2(_02096_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07365_ (.A1(net87),
    .A2(_02090_),
    .B(_02085_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07366_ (.A1(_02087_),
    .A2(_02097_),
    .B(_02098_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07367_ (.A1(\wb_counter[23] ),
    .A2(_02096_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07368_ (.A1(\wb_counter[24] ),
    .A2(_02099_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07369_ (.I(_02068_),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07370_ (.A1(net88),
    .A2(_02090_),
    .B(_02101_),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07371_ (.A1(_02087_),
    .A2(_02100_),
    .B(_02102_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07372_ (.I(_02000_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07373_ (.A1(\wb_counter[23] ),
    .A2(\wb_counter[24] ),
    .A3(_02096_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07374_ (.A1(\wb_counter[25] ),
    .A2(_02104_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07375_ (.I(_02018_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07376_ (.A1(net89),
    .A2(_02106_),
    .B(_02101_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07377_ (.A1(_02103_),
    .A2(_02105_),
    .B(_02107_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07378_ (.I(\wb_counter[25] ),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07379_ (.A1(_02108_),
    .A2(_02104_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07380_ (.A1(\wb_counter[26] ),
    .A2(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07381_ (.A1(net90),
    .A2(_02106_),
    .B(_02101_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07382_ (.A1(_02103_),
    .A2(_02110_),
    .B(_02111_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07383_ (.A1(\wb_counter[26] ),
    .A2(_02109_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07384_ (.A1(\wb_counter[27] ),
    .A2(_02112_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07385_ (.A1(net91),
    .A2(_02106_),
    .B(_02101_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07386_ (.A1(_02103_),
    .A2(_02113_),
    .B(_02114_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07387_ (.A1(\wb_counter[26] ),
    .A2(\wb_counter[27] ),
    .A3(_02109_),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07388_ (.A1(\wb_counter[28] ),
    .A2(_02115_),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07389_ (.I(_02068_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07390_ (.A1(net92),
    .A2(_02106_),
    .B(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07391_ (.A1(_02103_),
    .A2(_02116_),
    .B(net411),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07392_ (.I(\wb_counter[28] ),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07393_ (.A1(_02119_),
    .A2(_02115_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07394_ (.A1(\wb_counter[29] ),
    .A2(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07395_ (.A1(net93),
    .A2(_02019_),
    .B(_02117_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07396_ (.A1(_02011_),
    .A2(_02121_),
    .B(_02122_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07397_ (.A1(\wb_counter[29] ),
    .A2(_02120_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07398_ (.A1(\wb_counter[30] ),
    .A2(_02123_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07399_ (.A1(net95),
    .A2(_02019_),
    .B(_02117_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07400_ (.A1(_02011_),
    .A2(_02124_),
    .B(net405),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07401_ (.A1(\wb_counter[29] ),
    .A2(\wb_counter[30] ),
    .A3(_02120_),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07402_ (.A1(\wb_counter[31] ),
    .A2(_02126_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07403_ (.A1(net96),
    .A2(_02019_),
    .B(_02117_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07404_ (.A1(_02011_),
    .A2(_02127_),
    .B(_02128_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07405_ (.I(_01068_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07406_ (.A1(net240),
    .A2(_02129_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07407_ (.I(_01561_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07408_ (.A1(net221),
    .A2(_02131_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07409_ (.A1(_02130_),
    .A2(_02132_),
    .B(_01662_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07410_ (.A1(net247),
    .A2(net238),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07411_ (.I(_01066_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07412_ (.A1(net228),
    .A2(_02134_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07413_ (.A1(_01444_),
    .A2(_02133_),
    .A3(_02135_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07414_ (.A1(net248),
    .A2(_02129_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07415_ (.A1(net229),
    .A2(_02131_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07416_ (.A1(_02136_),
    .A2(_02137_),
    .B(_01662_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07417_ (.I(_01442_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07418_ (.I(_02138_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07419_ (.A1(net249),
    .A2(net238),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07420_ (.A1(net230),
    .A2(_02134_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07421_ (.A1(_02139_),
    .A2(_02140_),
    .A3(_02141_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07422_ (.A1(net250),
    .A2(_02129_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07423_ (.A1(net231),
    .A2(_02131_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07424_ (.A1(_02142_),
    .A2(_02143_),
    .B(_01662_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07425_ (.A1(net251),
    .A2(_02129_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07426_ (.A1(net232),
    .A2(_02134_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07427_ (.A1(_02139_),
    .A2(_02144_),
    .A3(_02145_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07428_ (.A1(net252),
    .A2(_01573_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07429_ (.A1(net233),
    .A2(_01562_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07430_ (.I(_01661_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07431_ (.A1(_02146_),
    .A2(_02147_),
    .B(_02148_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07432_ (.I(_02138_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07433_ (.A1(net234),
    .A2(_02131_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07434_ (.A1(_01026_),
    .A2(_02134_),
    .B(_02149_),
    .C(_02150_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07435_ (.A1(_01387_),
    .A2(_01660_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07436_ (.I(_01265_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07437_ (.I(_01237_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07438_ (.A1(_02153_),
    .A2(_01426_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07439_ (.I(_02154_),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07440_ (.I(_01228_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07441_ (.A1(_01424_),
    .A2(_02156_),
    .A3(_01374_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07442_ (.A1(_02155_),
    .A2(_02157_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07443_ (.A1(_02152_),
    .A2(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07444_ (.I(_02159_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07445_ (.A1(_01208_),
    .A2(_01145_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07446_ (.A1(_02161_),
    .A2(_01368_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07447_ (.I(_01264_),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07448_ (.I(_01288_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07449_ (.A1(_02163_),
    .A2(_02164_),
    .A3(_01227_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07450_ (.A1(_02162_),
    .A2(_02165_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07451_ (.A1(_01225_),
    .A2(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07452_ (.I(_02167_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07453_ (.I(_02168_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(_01204_),
    .A2(_01195_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07455_ (.I(_02170_),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07456_ (.A1(_02160_),
    .A2(_02169_),
    .B(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07457_ (.I(_01150_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07458_ (.I(_02159_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07459_ (.I(_01839_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07460_ (.I(_02175_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07461_ (.I(_02176_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07462_ (.A1(\as2650.debug_psu[0] ),
    .A2(\as2650.debug_psu[1] ),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07463_ (.I(_02178_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07464_ (.A1(_01835_),
    .A2(_01852_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07465_ (.A1(_02179_),
    .A2(_02180_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07466_ (.I(_02181_),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07467_ (.I(_02182_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07468_ (.I(_02183_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07469_ (.I(_02184_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07470_ (.I(_02185_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07471_ (.I(_02186_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07472_ (.I(_01838_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07473_ (.I(_02188_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07474_ (.I(_02189_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07475_ (.I(_02190_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07476_ (.I(\as2650.stack[0][13] ),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07477_ (.A1(_02191_),
    .A2(_02192_),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07478_ (.A1(_02177_),
    .A2(\as2650.stack[1][13] ),
    .B(_02187_),
    .C(_02193_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07479_ (.I(_02179_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07480_ (.I(_02195_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07481_ (.I(_02196_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07482_ (.I(_02197_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07483_ (.I(_02198_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07484_ (.I(_02199_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07485_ (.I(_02180_),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07486_ (.I(_02201_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07487_ (.I(_02202_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07488_ (.I(_02203_),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07489_ (.I(_02204_),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07490_ (.I(_02205_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07491_ (.A1(\as2650.debug_psu[2] ),
    .A2(_02178_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07492_ (.I(_02207_),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07493_ (.I(_02208_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07494_ (.I(_02209_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07495_ (.I(_02210_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07496_ (.I(_02211_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07497_ (.A1(\as2650.stack[3][13] ),
    .A2(_02200_),
    .B1(_02206_),
    .B2(\as2650.stack[2][13] ),
    .C(_02212_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07498_ (.I(\as2650.stack[4][13] ),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07499_ (.A1(_02191_),
    .A2(_02214_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07500_ (.A1(_02177_),
    .A2(\as2650.stack[5][13] ),
    .B(_02187_),
    .C(_02215_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07501_ (.I(_01861_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07502_ (.A1(_02217_),
    .A2(_02178_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07503_ (.I(_02218_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07504_ (.I(_02219_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07505_ (.I(_02220_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07506_ (.I(_02221_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07507_ (.I(_02222_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07508_ (.A1(\as2650.stack[7][13] ),
    .A2(_02200_),
    .B1(_02206_),
    .B2(\as2650.stack[6][13] ),
    .C(_02223_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07509_ (.A1(_02194_),
    .A2(_02213_),
    .B1(_02216_),
    .B2(_02224_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07510_ (.I(\as2650.stack[8][13] ),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07511_ (.A1(_02191_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07512_ (.A1(_02177_),
    .A2(\as2650.stack[9][13] ),
    .B(_02187_),
    .C(_02227_),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07513_ (.I(_02198_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07514_ (.I(_02229_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07515_ (.A1(\as2650.stack[11][13] ),
    .A2(_02230_),
    .B1(_02206_),
    .B2(\as2650.stack[10][13] ),
    .C(_02212_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07516_ (.I(_02190_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07517_ (.I(_01835_),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07518_ (.I(_02233_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07519_ (.I(_02234_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07520_ (.I(_02235_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07521_ (.I(_02236_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07522_ (.I(_02237_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07523_ (.I(_02238_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07524_ (.I(\as2650.stack[12][13] ),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07525_ (.A1(_02239_),
    .A2(_02240_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07526_ (.A1(_02232_),
    .A2(\as2650.stack[13][13] ),
    .B(_02187_),
    .C(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07527_ (.I(_02220_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07528_ (.I(_02243_),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07529_ (.A1(\as2650.stack[15][13] ),
    .A2(_02200_),
    .B1(_02206_),
    .B2(\as2650.stack[14][13] ),
    .C(_02244_),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07530_ (.A1(_02228_),
    .A2(_02231_),
    .B1(_02242_),
    .B2(_02245_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07531_ (.A1(_01861_),
    .A2(\as2650.debug_psu[3] ),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07532_ (.A1(_02179_),
    .A2(_02247_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07533_ (.A1(_01835_),
    .A2(_01852_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07534_ (.A1(_01861_),
    .A2(_02249_),
    .B(_01870_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07535_ (.A1(_02248_),
    .A2(_02250_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07536_ (.I(_02251_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07537_ (.I(_02252_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07538_ (.I(_02253_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07539_ (.I(_02254_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _07540_ (.I0(_02225_),
    .I1(_02246_),
    .S(_02255_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07541_ (.I(_00589_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07542_ (.A1(_02257_),
    .A2(_01188_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07543_ (.A1(_02258_),
    .A2(_01369_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07544_ (.I(_02259_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07545_ (.I(_02260_),
    .Z(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07546_ (.A1(_01421_),
    .A2(_02261_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07547_ (.A1(net216),
    .A2(_02174_),
    .B1(_02169_),
    .B2(_02256_),
    .C(_02262_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07548_ (.A1(_02173_),
    .A2(_02263_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07549_ (.A1(_01887_),
    .A2(_02172_),
    .B(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07550_ (.I(_01653_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07551_ (.I(_02164_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07552_ (.I(_02267_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07553_ (.I(_02268_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07554_ (.I(_01251_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07555_ (.A1(_02270_),
    .A2(_01452_),
    .A3(_01397_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07556_ (.A1(_01127_),
    .A2(_02153_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07557_ (.A1(_02271_),
    .A2(_02272_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07558_ (.A1(_02269_),
    .A2(_02273_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07559_ (.A1(_01399_),
    .A2(_02266_),
    .A3(_02274_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07560_ (.I(_02275_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07561_ (.A1(_02265_),
    .A2(_02276_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07562_ (.I(_01154_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07563_ (.I(_02278_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07564_ (.A1(_02279_),
    .A2(_01132_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07565_ (.A1(net63),
    .A2(_02279_),
    .B(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07566_ (.I(_02281_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07567_ (.I(_02152_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07568_ (.I(_02283_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07569_ (.I(_01126_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07570_ (.I(_02285_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07571_ (.I(_01237_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07572_ (.A1(_02286_),
    .A2(_02287_),
    .A3(_01422_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07573_ (.I(_02288_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07574_ (.A1(_02284_),
    .A2(_02289_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07575_ (.I(_02163_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07576_ (.A1(_02291_),
    .A2(_02282_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07577_ (.A1(_01887_),
    .A2(_02282_),
    .B(_02290_),
    .C(_02292_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07578_ (.I(_01411_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07579_ (.A1(_01168_),
    .A2(_02265_),
    .B(_02293_),
    .C(_02294_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07580_ (.A1(_02277_),
    .A2(_02295_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07581_ (.A1(_02151_),
    .A2(_02296_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07582_ (.I(_01201_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07583_ (.I(_02170_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07584_ (.I(_02298_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07585_ (.I(_02299_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07586_ (.I(_01532_),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07587_ (.I(_01086_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07588_ (.I(_02302_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07589_ (.I(_02303_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07590_ (.I(_01388_),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07591_ (.A1(\as2650.insin[0] ),
    .A2(_02300_),
    .B1(_02301_),
    .B2(_02304_),
    .C(_02305_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07592_ (.A1(_02297_),
    .A2(_02306_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07593_ (.I(_00860_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07594_ (.I(_02307_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07595_ (.I(_02308_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07596_ (.I(_02309_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07597_ (.A1(\as2650.insin[1] ),
    .A2(_02300_),
    .B1(_02301_),
    .B2(_02310_),
    .C(_02305_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07598_ (.A1(_02297_),
    .A2(_02311_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07599_ (.I(\as2650.is_interrupt_cycle ),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07600_ (.I(_02312_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07601_ (.I(_02313_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07602_ (.I(_01149_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07603_ (.I(_02315_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07604_ (.I(_02316_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07605_ (.I(_02315_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07606_ (.A1(_02318_),
    .A2(_01241_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _07607_ (.I0(net60),
    .I1(_01093_),
    .S(_01154_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07608_ (.I(_02320_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07609_ (.I(_02321_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07610_ (.I(_02322_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07611_ (.I(_02323_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07612_ (.A1(\as2650.insin[2] ),
    .A2(_02317_),
    .B1(_02319_),
    .B2(_02324_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07613_ (.A1(_02314_),
    .A2(_02325_),
    .B(_02148_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07614_ (.I(_01091_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07615_ (.I(_02326_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07616_ (.I(_02327_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07617_ (.I(_02328_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07618_ (.I(_02329_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07619_ (.A1(\as2650.insin[3] ),
    .A2(_02317_),
    .B1(_02319_),
    .B2(_02330_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07620_ (.A1(_02314_),
    .A2(_02331_),
    .B(_02148_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07621_ (.I(_01660_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07622_ (.I(_02332_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07623_ (.I(_02170_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07624_ (.I(_02334_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07625_ (.I(_01142_),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07626_ (.I(_02336_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07627_ (.I(_02337_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07628_ (.A1(\as2650.insin[4] ),
    .A2(_02335_),
    .B1(_02301_),
    .B2(_02338_),
    .C(_02305_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07629_ (.A1(_02333_),
    .A2(_02339_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07630_ (.I(_01134_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07631_ (.I(_02340_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07632_ (.I(_02341_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07633_ (.I(_02342_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07634_ (.A1(\as2650.insin[5] ),
    .A2(_02335_),
    .B1(_02301_),
    .B2(_02343_),
    .C(_01389_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07635_ (.A1(_02333_),
    .A2(_02344_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07636_ (.A1(_00678_),
    .A2(_00679_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07637_ (.I(_02345_),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07638_ (.I(_02346_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07639_ (.I(_01172_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07640_ (.A1(_01165_),
    .A2(_01416_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07641_ (.I(\as2650.PC[0] ),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07642_ (.I(_02350_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07643_ (.I(_02303_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07644_ (.A1(_02351_),
    .A2(_02352_),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07645_ (.A1(_01427_),
    .A2(_01267_),
    .A3(_01405_),
    .A4(_01374_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07646_ (.I(_02354_),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07647_ (.I(_02355_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07648_ (.I(_02356_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07649_ (.A1(_02350_),
    .A2(_02345_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07650_ (.A1(_02357_),
    .A2(_02358_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07651_ (.I(_02351_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07652_ (.A1(_02360_),
    .A2(_01376_),
    .B(_02346_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07653_ (.A1(_02359_),
    .A2(_02361_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07654_ (.I(_01409_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07655_ (.A1(_01657_),
    .A2(_02353_),
    .B1(_02362_),
    .B2(_02363_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07656_ (.A1(_01408_),
    .A2(_01656_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07657_ (.A1(_02349_),
    .A2(_02365_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07658_ (.A1(_02348_),
    .A2(_02349_),
    .A3(_02364_),
    .B1(_02366_),
    .B2(_00636_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07659_ (.I(_01393_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07660_ (.A1(_00636_),
    .A2(_02294_),
    .B(_02151_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07661_ (.A1(_02347_),
    .A2(_01395_),
    .B1(_02367_),
    .B2(_02368_),
    .C(_02369_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07662_ (.A1(_00981_),
    .A2(_01178_),
    .A3(_01457_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07663_ (.I(_02370_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07664_ (.I(_02371_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07665_ (.I(_01267_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07666_ (.A1(_02373_),
    .A2(_01258_),
    .A3(_01535_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07667_ (.A1(_02372_),
    .A2(_02374_),
    .B(\as2650.cpu_hidden_rom_enable ),
    .C(_01443_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07668_ (.A1(_01975_),
    .A2(_02139_),
    .B(_02375_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07669_ (.I(_01080_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07670_ (.I(_01392_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07671_ (.A1(_02377_),
    .A2(_02366_),
    .B(_01195_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07672_ (.I(_02378_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07673_ (.I(_00669_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07674_ (.I(_02380_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07675_ (.I(_01393_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07676_ (.I(_02382_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07677_ (.I(_01656_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07678_ (.A1(\as2650.PC[0] ),
    .A2(\as2650.PC[1] ),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07679_ (.I(_02385_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07680_ (.A1(_02308_),
    .A2(_02358_),
    .A3(_02386_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07681_ (.I(_02355_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07682_ (.I(_02355_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07683_ (.A1(_02389_),
    .A2(_02387_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07684_ (.A1(_02381_),
    .A2(_02388_),
    .B(_02390_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07685_ (.I(_01408_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07686_ (.A1(_02384_),
    .A2(_02387_),
    .B1(_02391_),
    .B2(_02392_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07687_ (.A1(_01165_),
    .A2(_01416_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07688_ (.A1(_01393_),
    .A2(_02394_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07689_ (.I(_02395_),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07690_ (.A1(_02381_),
    .A2(_02383_),
    .B1(_02393_),
    .B2(_02396_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07691_ (.I(_01387_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07692_ (.A1(\as2650.indirect_target[1] ),
    .A2(_02379_),
    .B1(_02397_),
    .B2(_02294_),
    .C(_02398_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07693_ (.I(\as2650.irqs_latch[6] ),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07694_ (.I(\as2650.irqs_latch[2] ),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07695_ (.A1(\as2650.irqs_latch[1] ),
    .A2(_02401_),
    .B(\as2650.irqs_latch[3] ),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07696_ (.I(\as2650.irqs_latch[5] ),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07697_ (.A1(\as2650.irqs_latch[4] ),
    .A2(_02402_),
    .B(_02403_),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07698_ (.A1(_02312_),
    .A2(\as2650.irqs_latch[7] ),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07699_ (.A1(_02400_),
    .A2(_02404_),
    .B(_02405_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07700_ (.A1(_02376_),
    .A2(_02399_),
    .A3(_02406_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07701_ (.I(_02378_),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07702_ (.I(_01095_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07703_ (.I(_02408_),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07704_ (.I(\as2650.PC[2] ),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07705_ (.A1(\as2650.PC[0] ),
    .A2(\as2650.PC[1] ),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07706_ (.A1(_02410_),
    .A2(_02411_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07707_ (.I(_02412_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07708_ (.A1(_00860_),
    .A2(_02385_),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07709_ (.A1(_02307_),
    .A2(_02385_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07710_ (.A1(_02358_),
    .A2(_02414_),
    .B(_02415_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07711_ (.A1(_01095_),
    .A2(_02413_),
    .A3(_02416_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07712_ (.A1(_02389_),
    .A2(_02417_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07713_ (.A1(_02408_),
    .A2(_02388_),
    .B(_02418_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07714_ (.A1(_01657_),
    .A2(_02417_),
    .B1(_02419_),
    .B2(_02363_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _07715_ (.A1(_02409_),
    .A2(_02383_),
    .B1(_02396_),
    .B2(_02420_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07716_ (.I(_01196_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07717_ (.A1(\as2650.indirect_target[2] ),
    .A2(_02407_),
    .B1(_02421_),
    .B2(_02422_),
    .C(_02398_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07718_ (.I(\as2650.irqs_latch[3] ),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07719_ (.A1(_02401_),
    .A2(_02424_),
    .B(\as2650.irqs_latch[4] ),
    .C(\as2650.irqs_latch[5] ),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07720_ (.A1(\as2650.irqs_latch[6] ),
    .A2(_02405_),
    .A3(_02425_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07721_ (.A1(_02376_),
    .A2(_02423_),
    .A3(_02426_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07722_ (.I(_02378_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07723_ (.I(_02395_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07724_ (.I(\as2650.PC[3] ),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07725_ (.I(\as2650.PC[1] ),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07726_ (.A1(_02350_),
    .A2(_02430_),
    .A3(_02410_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07727_ (.A1(_02429_),
    .A2(_02431_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07728_ (.I(_02432_),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07729_ (.A1(_02321_),
    .A2(_02412_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07730_ (.I(_02416_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07731_ (.A1(_02320_),
    .A2(_02412_),
    .B(_02435_),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07732_ (.A1(_02434_),
    .A2(_02436_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07733_ (.A1(_02327_),
    .A2(_02433_),
    .A3(_02437_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07734_ (.A1(_02356_),
    .A2(_02438_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07735_ (.A1(_02328_),
    .A2(_02388_),
    .B(_02439_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07736_ (.A1(_02384_),
    .A2(_02438_),
    .B1(_02440_),
    .B2(_01409_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07737_ (.A1(_02329_),
    .A2(_02382_),
    .B1(_02428_),
    .B2(_02441_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07738_ (.A1(_00629_),
    .A2(_02427_),
    .B1(_02442_),
    .B2(_01197_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07739_ (.A1(_02305_),
    .A2(_02443_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _07740_ (.A1(\as2650.irqs_latch[4] ),
    .A2(\as2650.irqs_latch[5] ),
    .A3(\as2650.irqs_latch[6] ),
    .A4(_02405_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07741_ (.A1(_02376_),
    .A2(_02444_),
    .A3(_02445_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07742_ (.A1(_01154_),
    .A2(_01140_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07743_ (.A1(net62),
    .A2(_02278_),
    .B(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07744_ (.I(_02447_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07745_ (.I(_02448_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07746_ (.I(_02449_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07747_ (.I(\as2650.PC[4] ),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07748_ (.A1(_00632_),
    .A2(_02431_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07749_ (.A1(_02451_),
    .A2(_02452_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07750_ (.I(_02432_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07751_ (.A1(_01156_),
    .A2(_02432_),
    .B1(_02436_),
    .B2(_02434_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07752_ (.A1(_01091_),
    .A2(_02454_),
    .B(_02455_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07753_ (.A1(_02448_),
    .A2(_02453_),
    .A3(_02456_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07754_ (.A1(_02389_),
    .A2(_02457_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07755_ (.A1(_02449_),
    .A2(_02357_),
    .B(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07756_ (.A1(_01657_),
    .A2(_02457_),
    .B1(_02459_),
    .B2(_02363_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07757_ (.A1(_02450_),
    .A2(_02383_),
    .B1(_02396_),
    .B2(_02460_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07758_ (.A1(\as2650.indirect_target[4] ),
    .A2(_02379_),
    .B1(_02461_),
    .B2(_01448_),
    .C(_01389_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07759_ (.A1(\as2650.ivectors_base[0] ),
    .A2(_02314_),
    .B(_01509_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07760_ (.A1(_02462_),
    .A2(_02463_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07761_ (.I(_01387_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07762_ (.I(_02464_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07763_ (.I(\as2650.indirect_target[5] ),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07764_ (.I(_02382_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07765_ (.I(\as2650.PC[5] ),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07766_ (.A1(_02451_),
    .A2(_02452_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _07767_ (.A1(_02468_),
    .A2(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07768_ (.I(\as2650.PC[4] ),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07769_ (.A1(_02471_),
    .A2(_02452_),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07770_ (.A1(_02447_),
    .A2(_02472_),
    .B(_02456_),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07771_ (.A1(_02336_),
    .A2(_02453_),
    .B(_02473_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07772_ (.A1(_02341_),
    .A2(_02470_),
    .A3(_02474_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07773_ (.A1(_02356_),
    .A2(_02475_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07774_ (.A1(_02342_),
    .A2(_02389_),
    .B(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07775_ (.A1(_02384_),
    .A2(_02475_),
    .B1(_02477_),
    .B2(_02392_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07776_ (.A1(_02343_),
    .A2(_02467_),
    .B1(_02396_),
    .B2(_02478_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07777_ (.A1(_02466_),
    .A2(_02407_),
    .B1(_02479_),
    .B2(_02422_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07778_ (.A1(_02465_),
    .A2(_02480_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07779_ (.I(_01508_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07780_ (.A1(\as2650.ivectors_base[1] ),
    .A2(_02314_),
    .B(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07781_ (.A1(_02481_),
    .A2(_02483_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07782_ (.I(_01121_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07783_ (.I(_02484_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07784_ (.I(_02485_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07785_ (.I(_02486_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07786_ (.I(_02487_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07787_ (.A1(_02278_),
    .A2(_01119_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07788_ (.A1(net64),
    .A2(_02278_),
    .B(_02489_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07789_ (.A1(\as2650.PC[4] ),
    .A2(_02468_),
    .A3(_02452_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07790_ (.A1(\as2650.PC[6] ),
    .A2(_02491_),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07791_ (.A1(_02490_),
    .A2(_02492_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07792_ (.A1(_02468_),
    .A2(_02469_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07793_ (.A1(_02281_),
    .A2(_02494_),
    .B(_02474_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07794_ (.A1(_02340_),
    .A2(_02470_),
    .B(_02495_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07795_ (.A1(_02493_),
    .A2(_02496_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07796_ (.A1(_01376_),
    .A2(_02365_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07797_ (.A1(_02487_),
    .A2(_02354_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07798_ (.I(_02499_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07799_ (.A1(_02497_),
    .A2(_02498_),
    .B1(_02500_),
    .B2(_02392_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07800_ (.A1(_02488_),
    .A2(_02467_),
    .B1(_02428_),
    .B2(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07801_ (.A1(_00623_),
    .A2(_02407_),
    .B1(_02502_),
    .B2(_02422_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07802_ (.A1(_02465_),
    .A2(_02503_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07803_ (.I(_02312_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07804_ (.A1(\as2650.ivectors_base[2] ),
    .A2(_02505_),
    .B(_02482_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07805_ (.A1(_02504_),
    .A2(_02506_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07806_ (.I(\as2650.indirect_target[7] ),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07807_ (.I(_01403_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07808_ (.I(_02508_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07809_ (.I(\as2650.PC[6] ),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07810_ (.A1(_02510_),
    .A2(\as2650.PC[7] ),
    .A3(_02491_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07811_ (.A1(_02510_),
    .A2(_02491_),
    .B(\as2650.PC[7] ),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07812_ (.A1(_02511_),
    .A2(_02512_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07813_ (.I(_02513_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07814_ (.A1(_02493_),
    .A2(_02496_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07815_ (.A1(_02484_),
    .A2(_02492_),
    .B(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07816_ (.A1(_02486_),
    .A2(_02514_),
    .A3(_02516_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07817_ (.A1(_02356_),
    .A2(_02517_),
    .B(_02500_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07818_ (.I(_02518_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07819_ (.A1(_02384_),
    .A2(_02517_),
    .B1(_02519_),
    .B2(_01409_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07820_ (.A1(_02509_),
    .A2(_02467_),
    .B1(_02428_),
    .B2(_02520_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07821_ (.I(_01196_),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07822_ (.A1(_02507_),
    .A2(_02427_),
    .B1(_02521_),
    .B2(_02522_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07823_ (.A1(_02465_),
    .A2(_02523_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07824_ (.A1(\as2650.ivectors_base[3] ),
    .A2(_02505_),
    .B(_02482_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07825_ (.A1(_02524_),
    .A2(_02525_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07826_ (.I(\as2650.indirect_target[8] ),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07827_ (.I(_02490_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07828_ (.I(\as2650.PC[8] ),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07829_ (.A1(_02528_),
    .A2(_02511_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07830_ (.A1(_02527_),
    .A2(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07831_ (.A1(_02527_),
    .A2(_02513_),
    .B(_02516_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07832_ (.A1(_02485_),
    .A2(_02514_),
    .B(_02531_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07833_ (.A1(_02530_),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07834_ (.A1(_02392_),
    .A2(_02500_),
    .B1(_02533_),
    .B2(_02498_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07835_ (.A1(\as2650.instruction_args_latch[8] ),
    .A2(_02467_),
    .B1(_02428_),
    .B2(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07836_ (.A1(_02526_),
    .A2(_02427_),
    .B1(_02535_),
    .B2(_02522_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07837_ (.A1(_02465_),
    .A2(_02536_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07838_ (.A1(\as2650.ivectors_base[4] ),
    .A2(_02505_),
    .B(_02482_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07839_ (.A1(_02537_),
    .A2(_02538_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07840_ (.I(\as2650.ivectors_base[5] ),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07841_ (.I(_02398_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07842_ (.I(\as2650.instruction_args_latch[9] ),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07843_ (.A1(_02541_),
    .A2(_01395_),
    .B(_02398_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07844_ (.I(\as2650.PC[9] ),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07845_ (.A1(_02528_),
    .A2(_02511_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07846_ (.A1(_02543_),
    .A2(_02544_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07847_ (.A1(_02527_),
    .A2(_02545_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07848_ (.I(_02529_),
    .Z(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07849_ (.A1(_02487_),
    .A2(_02547_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07850_ (.A1(_02548_),
    .A2(_02532_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07851_ (.A1(_02488_),
    .A2(_02547_),
    .B(_02549_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07852_ (.A1(_02546_),
    .A2(_02550_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07853_ (.I(_02498_),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07854_ (.A1(_02394_),
    .A2(_02552_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07855_ (.A1(_01488_),
    .A2(_02377_),
    .A3(_02553_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07856_ (.A1(\as2650.indirect_target[9] ),
    .A2(_02379_),
    .B1(_02551_),
    .B2(_02554_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07857_ (.A1(_02539_),
    .A2(_02540_),
    .B1(_02542_),
    .B2(_02555_),
    .C(_01081_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07858_ (.I(\as2650.ivectors_base[6] ),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07859_ (.I(_02527_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07860_ (.I(\as2650.PC[10] ),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07861_ (.A1(\as2650.PC[8] ),
    .A2(_02543_),
    .A3(_02511_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07862_ (.A1(_02558_),
    .A2(_02559_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07863_ (.A1(_02557_),
    .A2(_02560_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07864_ (.I(_02560_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07865_ (.A1(_02557_),
    .A2(_02562_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07866_ (.A1(_02561_),
    .A2(_02563_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07867_ (.A1(_02547_),
    .A2(_02545_),
    .B(_02485_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07868_ (.A1(_02530_),
    .A2(_02532_),
    .A3(_02546_),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07869_ (.A1(_02565_),
    .A2(_02566_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07870_ (.A1(_02564_),
    .A2(_02567_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07871_ (.A1(_02554_),
    .A2(_02568_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07872_ (.I(\as2650.instruction_args_latch[10] ),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07873_ (.A1(_02570_),
    .A2(_01395_),
    .B1(_02407_),
    .B2(\as2650.indirect_target[10] ),
    .C(_02464_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07874_ (.I(_01078_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07875_ (.I(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07876_ (.I(_02573_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07877_ (.A1(_02556_),
    .A2(_02540_),
    .B1(_02569_),
    .B2(_02571_),
    .C(_02574_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07878_ (.A1(_01411_),
    .A2(_02382_),
    .A3(_02394_),
    .A4(_02552_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07879_ (.I(\as2650.PC[11] ),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07880_ (.I(_02558_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07881_ (.A1(_02577_),
    .A2(_02559_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07882_ (.A1(_02576_),
    .A2(_02578_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07883_ (.A1(_02484_),
    .A2(_02579_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07884_ (.I(_02561_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07885_ (.A1(_02581_),
    .A2(_02567_),
    .B(_02563_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07886_ (.A1(_02580_),
    .A2(_02582_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07887_ (.A1(\as2650.indirect_target[11] ),
    .A2(_02427_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07888_ (.I(\as2650.instruction_args_latch[11] ),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07889_ (.I(_01394_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07890_ (.A1(_02585_),
    .A2(_02586_),
    .B(_01388_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07891_ (.A1(_02575_),
    .A2(_02583_),
    .B(_02584_),
    .C(_02587_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07892_ (.A1(\as2650.ivectors_base[7] ),
    .A2(_02505_),
    .B(_02588_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07893_ (.A1(_02333_),
    .A2(_02589_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07894_ (.I(_02557_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07895_ (.A1(_02590_),
    .A2(_02579_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07896_ (.A1(_02564_),
    .A2(_02580_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07897_ (.A1(_02566_),
    .A2(_02592_),
    .B(_02565_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07898_ (.A1(_02487_),
    .A2(_02593_),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07899_ (.A1(_02591_),
    .A2(_02593_),
    .B(_02594_),
    .C(_02561_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07900_ (.I(\as2650.PC[12] ),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07901_ (.A1(_02576_),
    .A2(_02578_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _07902_ (.A1(_02596_),
    .A2(_02597_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07903_ (.A1(_02595_),
    .A2(_02598_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07904_ (.I(\as2650.instruction_args_latch[12] ),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07905_ (.A1(_02600_),
    .A2(_02586_),
    .B1(_02378_),
    .B2(\as2650.indirect_target[12] ),
    .C(_01388_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07906_ (.A1(_02575_),
    .A2(_02599_),
    .B(_02601_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07907_ (.A1(\as2650.ivectors_base[8] ),
    .A2(_02313_),
    .B(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07908_ (.A1(_02333_),
    .A2(_02603_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07909_ (.I(\as2650.ivectors_base[9] ),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07910_ (.I(\as2650.indirect_target[13] ),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07911_ (.I(_02266_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07912_ (.A1(_00592_),
    .A2(_01417_),
    .A3(_02606_),
    .A4(_02552_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07913_ (.A1(_02605_),
    .A2(_02366_),
    .B(_02607_),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07914_ (.A1(_02368_),
    .A2(_02608_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07915_ (.I(_01172_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07916_ (.I(_02610_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07917_ (.I(\as2650.instruction_args_latch[13] ),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07918_ (.I(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07919_ (.I(_02613_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07920_ (.I(_01401_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07921_ (.A1(_00592_),
    .A2(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07922_ (.A1(_02614_),
    .A2(_02615_),
    .B(_02616_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07923_ (.A1(\as2650.indirect_target[13] ),
    .A2(_02611_),
    .B1(_02586_),
    .B2(_02617_),
    .C(_02464_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07924_ (.A1(_02604_),
    .A2(_02540_),
    .B1(_02609_),
    .B2(_02618_),
    .C(_02574_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07925_ (.I(\as2650.ivectors_base[10] ),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07926_ (.A1(\as2650.page_reg[1] ),
    .A2(_01417_),
    .A3(_02606_),
    .A4(_02552_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07927_ (.A1(_00930_),
    .A2(_02366_),
    .B(_02620_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07928_ (.A1(_02368_),
    .A2(_02621_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07929_ (.I(_00925_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07930_ (.A1(\as2650.page_reg[1] ),
    .A2(_02615_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07931_ (.A1(_02623_),
    .A2(_02615_),
    .B(_02624_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07932_ (.A1(\as2650.indirect_target[14] ),
    .A2(_02611_),
    .B1(_02586_),
    .B2(_02625_),
    .C(_02464_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07933_ (.A1(_02619_),
    .A2(_02540_),
    .B1(_02622_),
    .B2(_02626_),
    .C(_02574_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07934_ (.I(\as2650.page_reg[2] ),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07935_ (.A1(_02368_),
    .A2(_02553_),
    .B(_02627_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07936_ (.A1(\as2650.indirect_target[15] ),
    .A2(_02379_),
    .B1(_02628_),
    .B2(_02294_),
    .C(_01389_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07937_ (.I(_01550_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07938_ (.I(_02630_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07939_ (.A1(\as2650.ivectors_base[11] ),
    .A2(_02313_),
    .B(_02631_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07940_ (.A1(_02629_),
    .A2(_02632_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07941_ (.I(\as2650.instruction_args_latch[14] ),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07942_ (.A1(\as2650.instruction_args_latch[13] ),
    .A2(_02633_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07943_ (.A1(_01402_),
    .A2(_01169_),
    .A3(_01222_),
    .A4(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07944_ (.I(_02635_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07945_ (.A1(_01648_),
    .A2(\as2650.indexed_cyc[0] ),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07946_ (.A1(_02636_),
    .A2(_02637_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07947_ (.I(_02612_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07948_ (.I(_02639_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07949_ (.I(_02640_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07950_ (.A1(_02612_),
    .A2(_02633_),
    .B(_00940_),
    .C(_01401_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07951_ (.A1(_01230_),
    .A2(_01233_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07952_ (.I(_02643_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _07953_ (.A1(_02257_),
    .A2(_02644_),
    .A3(_01146_),
    .A4(_01427_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07954_ (.A1(_02642_),
    .A2(_02645_),
    .B(_01377_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07955_ (.A1(_02641_),
    .A2(_02636_),
    .A3(_02646_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07956_ (.I(_00650_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07957_ (.A1(_02648_),
    .A2(_02348_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07958_ (.I(_01080_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07959_ (.A1(_02638_),
    .A2(_02647_),
    .B(_02649_),
    .C(_02650_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07960_ (.A1(_01648_),
    .A2(\as2650.indexed_cyc[1] ),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07961_ (.A1(_02636_),
    .A2(_02651_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07962_ (.I(_02633_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07963_ (.A1(_02653_),
    .A2(_02636_),
    .A3(_02646_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07964_ (.A1(_02652_),
    .A2(_02654_),
    .B(_01081_),
    .C(_02649_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07965_ (.A1(_01167_),
    .A2(_01191_),
    .A3(_02363_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07966_ (.A1(_02383_),
    .A2(_02655_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07967_ (.A1(_01648_),
    .A2(_01402_),
    .B1(_02522_),
    .B2(_02656_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07968_ (.A1(_02649_),
    .A2(_02657_),
    .B(_02313_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07969_ (.A1(_01509_),
    .A2(_02658_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07970_ (.I(_02659_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07971_ (.I(_02270_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07972_ (.I(_02660_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07973_ (.A1(_01647_),
    .A2(_01250_),
    .B(_02661_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07974_ (.A1(_02335_),
    .A2(_01269_),
    .B(_02662_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07975_ (.A1(_01455_),
    .A2(_01458_),
    .A3(_02663_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07976_ (.A1(_02661_),
    .A2(_01505_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07977_ (.A1(_02664_),
    .A2(_02665_),
    .B(_02148_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07978_ (.I(_02332_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07979_ (.I(_01534_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07980_ (.I(_02667_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07981_ (.I(_02668_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07982_ (.A1(_01148_),
    .A2(_02669_),
    .B(net213),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07983_ (.A1(_02666_),
    .A2(_02670_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07984_ (.I(\as2650.warmup[1] ),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07985_ (.A1(\as2650.warmup[0] ),
    .A2(_02671_),
    .B(_01023_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07986_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07987_ (.A1(_01023_),
    .A2(_02672_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07988_ (.A1(_01205_),
    .A2(_01411_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07989_ (.I(_02673_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07990_ (.I(_02610_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07991_ (.A1(_01456_),
    .A2(_00735_),
    .A3(_01243_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07992_ (.A1(_01194_),
    .A2(_02304_),
    .B(_02676_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07993_ (.A1(_01204_),
    .A2(_01193_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07994_ (.I(_02678_),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07995_ (.A1(_01035_),
    .A2(_02679_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07996_ (.A1(_02675_),
    .A2(_02677_),
    .B(_02680_),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07997_ (.I(_00650_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07998_ (.A1(_01035_),
    .A2(_02674_),
    .B1(_02681_),
    .B2(_02682_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07999_ (.A1(_02666_),
    .A2(_02683_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08000_ (.I(_02673_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08001_ (.I(_01193_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08002_ (.A1(_02685_),
    .A2(_00753_),
    .A3(_01243_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08003_ (.A1(_01194_),
    .A2(_02310_),
    .B(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08004_ (.A1(\as2650.instruction_args_latch[1] ),
    .A2(_02679_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08005_ (.A1(_02675_),
    .A2(_02687_),
    .B(_02688_),
    .ZN(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08006_ (.A1(\as2650.instruction_args_latch[1] ),
    .A2(_02684_),
    .B1(_02689_),
    .B2(_02682_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08007_ (.A1(_02666_),
    .A2(_02690_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08008_ (.A1(_02685_),
    .A2(_00777_),
    .A3(_01243_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08009_ (.A1(_01194_),
    .A2(_02324_),
    .B(_02691_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08010_ (.A1(\as2650.instruction_args_latch[2] ),
    .A2(_02679_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08011_ (.A1(_02675_),
    .A2(_02692_),
    .B(_02693_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08012_ (.A1(\as2650.instruction_args_latch[2] ),
    .A2(_02684_),
    .B1(_02694_),
    .B2(_02682_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08013_ (.A1(_02666_),
    .A2(_02695_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08014_ (.I(_01660_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08015_ (.I(_02696_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08016_ (.I(_01242_),
    .Z(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08017_ (.A1(_02685_),
    .A2(_00800_),
    .A3(_02698_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08018_ (.A1(_01456_),
    .A2(_02330_),
    .B(_02699_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08019_ (.A1(\as2650.instruction_args_latch[3] ),
    .A2(_02679_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08020_ (.A1(_02675_),
    .A2(_02700_),
    .B(_02701_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08021_ (.A1(\as2650.instruction_args_latch[3] ),
    .A2(_02684_),
    .B1(_02702_),
    .B2(_02682_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08022_ (.A1(_02697_),
    .A2(_02703_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08023_ (.I(_02678_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _08024_ (.I(_00982_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08025_ (.I(_02705_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08026_ (.A1(_02706_),
    .A2(net200),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08027_ (.A1(_02706_),
    .A2(_02450_),
    .B1(_02698_),
    .B2(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08028_ (.A1(\as2650.instruction_args_latch[4] ),
    .A2(_02704_),
    .B1(_01197_),
    .B2(_02708_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08029_ (.A1(_01218_),
    .A2(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08030_ (.A1(\as2650.instruction_args_latch[4] ),
    .A2(_02674_),
    .B(_02710_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08031_ (.A1(_02697_),
    .A2(_02711_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08032_ (.I(_02610_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08033_ (.A1(_02685_),
    .A2(_00846_),
    .A3(_02698_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08034_ (.A1(_01456_),
    .A2(_02343_),
    .B(_02713_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08035_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_02704_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08036_ (.A1(_02712_),
    .A2(_02714_),
    .B(_02715_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08037_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_02684_),
    .B1(_02716_),
    .B2(_02648_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08038_ (.A1(_02697_),
    .A2(_02717_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _08039_ (.I(_02590_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08040_ (.I(_02718_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08041_ (.A1(_02705_),
    .A2(net202),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08042_ (.A1(_02706_),
    .A2(_02719_),
    .B1(_02698_),
    .B2(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08043_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_02704_),
    .B1(_01447_),
    .B2(_02721_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08044_ (.A1(_01218_),
    .A2(_02722_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08045_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_02674_),
    .B(_02723_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08046_ (.A1(_02697_),
    .A2(_02724_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08047_ (.I(_02696_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08048_ (.A1(_02279_),
    .A2(_01108_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08049_ (.A1(net65),
    .A2(_02279_),
    .B(_02726_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08050_ (.I(_02727_),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08051_ (.I(_02728_),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08052_ (.A1(_02705_),
    .A2(net203),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08053_ (.A1(_02706_),
    .A2(_02729_),
    .B1(_01242_),
    .B2(_02730_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08054_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_02704_),
    .B1(_01447_),
    .B2(_02731_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08055_ (.A1(_01218_),
    .A2(_02732_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08056_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_02674_),
    .B(_02733_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08057_ (.A1(_02725_),
    .A2(_02734_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08058_ (.I(_02648_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08059_ (.I(_01205_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08060_ (.I(_01165_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08061_ (.I(_02737_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08062_ (.I(_01166_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08063_ (.A1(_01166_),
    .A2(_01242_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08064_ (.I(_02740_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08065_ (.A1(_02739_),
    .A2(_02304_),
    .B1(net204),
    .B2(_02741_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08066_ (.A1(_02736_),
    .A2(_02738_),
    .A3(_00899_),
    .B1(_02712_),
    .B2(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08067_ (.A1(_02735_),
    .A2(_02743_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08068_ (.I(_01647_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08069_ (.I(_02745_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08070_ (.A1(_02746_),
    .A2(\as2650.instruction_args_latch[8] ),
    .A3(_01505_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08071_ (.I(_01661_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08072_ (.A1(_02744_),
    .A2(_02747_),
    .B(_02748_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08073_ (.I(_02541_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08074_ (.I(_02610_),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08075_ (.A1(_02739_),
    .A2(_02310_),
    .B1(net205),
    .B2(_02741_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08076_ (.A1(_02736_),
    .A2(_02738_),
    .A3(_02749_),
    .B1(_02750_),
    .B2(_02751_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08077_ (.A1(_02735_),
    .A2(_02752_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08078_ (.A1(_02746_),
    .A2(_02541_),
    .A3(_01505_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08079_ (.A1(_02753_),
    .A2(_02754_),
    .B(_02748_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08080_ (.A1(_02745_),
    .A2(_02570_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08081_ (.I(_01166_),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08082_ (.I(_02740_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08083_ (.A1(_02756_),
    .A2(_02324_),
    .B1(_02757_),
    .B2(net206),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08084_ (.A1(_01168_),
    .A2(_02755_),
    .B1(_02758_),
    .B2(_02712_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08085_ (.A1(_02735_),
    .A2(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08086_ (.I(_02348_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08087_ (.A1(_02746_),
    .A2(_02570_),
    .A3(_02761_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08088_ (.A1(_02760_),
    .A2(_02762_),
    .B(_02748_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08089_ (.A1(_02745_),
    .A2(_02585_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08090_ (.A1(_01167_),
    .A2(_02330_),
    .B1(_02757_),
    .B2(net207),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08091_ (.A1(_02738_),
    .A2(_02763_),
    .B1(_02764_),
    .B2(_02712_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08092_ (.A1(_02735_),
    .A2(_02765_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08093_ (.A1(_02746_),
    .A2(_02585_),
    .A3(_02761_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08094_ (.A1(_02766_),
    .A2(_02767_),
    .B(_02748_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08095_ (.I(_02648_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08096_ (.I(_02737_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08097_ (.I(_02600_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08098_ (.A1(_02739_),
    .A2(_02338_),
    .B1(_02741_),
    .B2(net208),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08099_ (.A1(_02736_),
    .A2(_02769_),
    .A3(_02770_),
    .B1(_02750_),
    .B2(_02771_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(_02768_),
    .A2(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08101_ (.I(_02745_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08102_ (.A1(_02774_),
    .A2(_02600_),
    .A3(_02761_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08103_ (.I(_01661_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08104_ (.A1(_02773_),
    .A2(_02775_),
    .B(_02776_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08105_ (.A1(_02756_),
    .A2(_02343_),
    .B1(_02741_),
    .B2(net209),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08106_ (.A1(_02736_),
    .A2(_02769_),
    .A3(_02614_),
    .B1(_02750_),
    .B2(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08107_ (.A1(_02768_),
    .A2(_02778_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08108_ (.A1(_02774_),
    .A2(_02641_),
    .A3(_02761_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08109_ (.A1(_02779_),
    .A2(_02780_),
    .B(_02776_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08110_ (.A1(_02756_),
    .A2(_02488_),
    .B1(_02757_),
    .B2(net211),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08111_ (.A1(_01206_),
    .A2(_02769_),
    .A3(_02623_),
    .B1(_02750_),
    .B2(_02781_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08112_ (.A1(_02768_),
    .A2(_02782_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08113_ (.A1(_02774_),
    .A2(_02653_),
    .A3(_02611_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08114_ (.A1(_02783_),
    .A2(_02784_),
    .B(_02776_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08115_ (.A1(_02756_),
    .A2(_02509_),
    .B1(_02757_),
    .B2(net212),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08116_ (.A1(_01206_),
    .A2(_02769_),
    .A3(_00939_),
    .B1(_02348_),
    .B2(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08117_ (.A1(_02768_),
    .A2(_02786_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08118_ (.A1(_02774_),
    .A2(\as2650.instruction_args_latch[15] ),
    .A3(_02611_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08119_ (.A1(_02787_),
    .A2(_02788_),
    .B(_02776_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08120_ (.A1(_01401_),
    .A2(_01223_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08121_ (.A1(_00981_),
    .A2(_01179_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08122_ (.A1(_02789_),
    .A2(_02790_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08123_ (.I(_02791_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08124_ (.I(_02792_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08125_ (.I(_01379_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08126_ (.I(_02794_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08127_ (.I(_02795_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08128_ (.A1(net212),
    .A2(_01403_),
    .A3(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08129_ (.A1(net211),
    .A2(_02795_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08130_ (.A1(_02557_),
    .A2(_02798_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08131_ (.A1(net209),
    .A2(_02340_),
    .A3(_02796_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08132_ (.A1(net208),
    .A2(_02794_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08133_ (.A1(_02448_),
    .A2(_02801_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08134_ (.A1(net207),
    .A2(_02326_),
    .A3(_02795_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08135_ (.A1(net206),
    .A2(_01378_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08136_ (.A1(_01095_),
    .A2(_02804_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08137_ (.A1(_02307_),
    .A2(net205),
    .A3(_02794_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08138_ (.A1(net205),
    .A2(_01378_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08139_ (.A1(_02380_),
    .A2(_02807_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08140_ (.A1(_02302_),
    .A2(_00739_),
    .A3(_01379_),
    .A4(_02808_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08141_ (.A1(_02321_),
    .A2(_02804_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08142_ (.A1(_02806_),
    .A2(_02809_),
    .B(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08143_ (.I(_01156_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08144_ (.A1(net207),
    .A2(_01379_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08145_ (.A1(_02812_),
    .A2(_02813_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08146_ (.A1(_02805_),
    .A2(_02811_),
    .B(_02814_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08147_ (.A1(_02336_),
    .A2(_02801_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08148_ (.A1(_02803_),
    .A2(_02815_),
    .B(_02816_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08149_ (.A1(net209),
    .A2(_02794_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08150_ (.A1(_02281_),
    .A2(_02818_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08151_ (.A1(_02802_),
    .A2(_02817_),
    .B(_02819_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08152_ (.A1(_02484_),
    .A2(_02798_),
    .Z(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08153_ (.A1(_02800_),
    .A2(_02820_),
    .B(_02821_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08154_ (.A1(net212),
    .A2(_02795_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08155_ (.A1(_02727_),
    .A2(_02823_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08156_ (.A1(_02799_),
    .A2(_02822_),
    .B(_02824_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08157_ (.A1(_02797_),
    .A2(_02825_),
    .B(_00899_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _08158_ (.A1(\as2650.instruction_args_latch[9] ),
    .A2(\as2650.instruction_args_latch[10] ),
    .A3(_02826_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08159_ (.A1(\as2650.instruction_args_latch[11] ),
    .A2(\as2650.instruction_args_latch[12] ),
    .A3(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08160_ (.A1(_02641_),
    .A2(_02828_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08161_ (.I(_00592_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08162_ (.I(_02260_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08163_ (.A1(_01150_),
    .A2(_02831_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08164_ (.A1(_01189_),
    .A2(_01454_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08165_ (.I(_02833_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08166_ (.I(_02834_),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08167_ (.A1(_02357_),
    .A2(_01650_),
    .A3(_02835_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08168_ (.A1(_02256_),
    .A2(_02832_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08169_ (.A1(_02830_),
    .A2(_02832_),
    .B(_02836_),
    .C(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08170_ (.A1(_02792_),
    .A2(_02838_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08171_ (.A1(_02793_),
    .A2(_02829_),
    .B(_02839_),
    .C(_02650_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08172_ (.I(_02371_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08173_ (.I(_02832_),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08174_ (.I(_02183_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08175_ (.I(_02842_),
    .Z(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08176_ (.I(_02843_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08177_ (.I(_02844_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08178_ (.I(_02845_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08179_ (.I(_02235_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08180_ (.I(_02847_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08181_ (.I(_02848_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08182_ (.I(_02849_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08183_ (.I(_02850_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08184_ (.I(\as2650.stack[0][14] ),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08185_ (.A1(_02851_),
    .A2(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08186_ (.A1(_01843_),
    .A2(\as2650.stack[1][14] ),
    .B(_02846_),
    .C(_02853_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08187_ (.I(_02196_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08188_ (.I(_02855_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08189_ (.I(_02856_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08190_ (.I(_02857_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08191_ (.I(_02858_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08192_ (.I(_02202_),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08193_ (.I(_02860_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08194_ (.I(_02861_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08195_ (.I(_02862_),
    .Z(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08196_ (.I(_02863_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08197_ (.I(_02210_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08198_ (.I(_02865_),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08199_ (.I(_02866_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08200_ (.A1(\as2650.stack[3][14] ),
    .A2(_02859_),
    .B1(_02864_),
    .B2(\as2650.stack[2][14] ),
    .C(_02867_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08201_ (.I(_01841_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08202_ (.I(_02869_),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08203_ (.I(_02845_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08204_ (.I(_02850_),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08205_ (.I(\as2650.stack[4][14] ),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08206_ (.A1(_02872_),
    .A2(_02873_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08207_ (.A1(_02870_),
    .A2(\as2650.stack[5][14] ),
    .B(_02871_),
    .C(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08208_ (.I(_02858_),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08209_ (.I(_02863_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08210_ (.I(_02244_),
    .Z(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08211_ (.A1(\as2650.stack[7][14] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\as2650.stack[6][14] ),
    .C(_02878_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08212_ (.A1(_02854_),
    .A2(_02868_),
    .B1(_02875_),
    .B2(_02879_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08213_ (.I(\as2650.stack[8][14] ),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08214_ (.A1(_02851_),
    .A2(_02881_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08215_ (.A1(_02870_),
    .A2(\as2650.stack[9][14] ),
    .B(_02846_),
    .C(_02882_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08216_ (.A1(\as2650.stack[11][14] ),
    .A2(_02859_),
    .B1(_02864_),
    .B2(\as2650.stack[10][14] ),
    .C(_02867_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08217_ (.I(_01841_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08218_ (.I(_02885_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08219_ (.I(\as2650.stack[12][14] ),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08220_ (.A1(_02872_),
    .A2(_02887_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08221_ (.A1(_02886_),
    .A2(\as2650.stack[13][14] ),
    .B(_02871_),
    .C(_02888_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08222_ (.A1(\as2650.stack[15][14] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\as2650.stack[14][14] ),
    .C(_02878_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08223_ (.A1(_02883_),
    .A2(_02884_),
    .B1(_02889_),
    .B2(_02890_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08224_ (.I(_02255_),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08225_ (.I0(_02880_),
    .I1(_02891_),
    .S(_02892_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08226_ (.A1(_00932_),
    .A2(_02841_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08227_ (.I(_02836_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08228_ (.A1(_02841_),
    .A2(_02893_),
    .B(_02894_),
    .C(_02895_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08229_ (.I(_02828_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08230_ (.A1(_02641_),
    .A2(_02653_),
    .A3(_02897_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08231_ (.A1(_02614_),
    .A2(_02828_),
    .B(_02623_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08232_ (.A1(_02898_),
    .A2(_02899_),
    .B(_02371_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08233_ (.I(_01201_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08234_ (.A1(_02840_),
    .A2(_02896_),
    .B(_02900_),
    .C(_02901_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08235_ (.I(\as2650.stack[0][15] ),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08236_ (.A1(_02851_),
    .A2(_02902_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08237_ (.A1(_02870_),
    .A2(\as2650.stack[1][15] ),
    .B(_02846_),
    .C(_02903_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08238_ (.A1(\as2650.stack[3][15] ),
    .A2(_02859_),
    .B1(_02864_),
    .B2(\as2650.stack[2][15] ),
    .C(_02867_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08239_ (.I(\as2650.stack[4][15] ),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08240_ (.A1(_02872_),
    .A2(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08241_ (.A1(_02886_),
    .A2(\as2650.stack[5][15] ),
    .B(_02871_),
    .C(_02907_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08242_ (.A1(\as2650.stack[7][15] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\as2650.stack[6][15] ),
    .C(_02878_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08243_ (.A1(_02904_),
    .A2(_02905_),
    .B1(_02908_),
    .B2(_02909_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08244_ (.I(\as2650.stack[8][15] ),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08245_ (.A1(_02872_),
    .A2(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08246_ (.A1(_02870_),
    .A2(\as2650.stack[9][15] ),
    .B(_02846_),
    .C(_02912_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08247_ (.I(_02198_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08248_ (.I(_02914_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08249_ (.A1(\as2650.stack[11][15] ),
    .A2(_02915_),
    .B1(_02864_),
    .B2(\as2650.stack[10][15] ),
    .C(_02867_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08250_ (.I(_02849_),
    .Z(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08251_ (.I(_02917_),
    .Z(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08252_ (.I(\as2650.stack[12][15] ),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08253_ (.A1(_02918_),
    .A2(_02919_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08254_ (.A1(_02886_),
    .A2(\as2650.stack[13][15] ),
    .B(_02871_),
    .C(_02920_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08255_ (.A1(\as2650.stack[15][15] ),
    .A2(_02859_),
    .B1(_02877_),
    .B2(\as2650.stack[14][15] ),
    .C(_02223_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08256_ (.A1(_02913_),
    .A2(_02916_),
    .B1(_02921_),
    .B2(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08257_ (.I0(_02910_),
    .I1(_02923_),
    .S(_02892_),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08258_ (.A1(_02627_),
    .A2(_02841_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08259_ (.A1(_02841_),
    .A2(_02924_),
    .B(_02925_),
    .C(_02895_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08260_ (.I(_00942_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08261_ (.A1(_02927_),
    .A2(_02898_),
    .Z(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08262_ (.A1(_02372_),
    .A2(_02928_),
    .B(_02631_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08263_ (.A1(_02840_),
    .A2(_02926_),
    .B(_02929_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08264_ (.I(_02156_),
    .Z(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08265_ (.A1(_02661_),
    .A2(_02930_),
    .A3(_01240_),
    .A4(_02373_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08266_ (.A1(_01426_),
    .A2(_02161_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08267_ (.I(_02152_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08268_ (.A1(_02660_),
    .A2(_01424_),
    .A3(_02933_),
    .A4(_02930_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08269_ (.A1(_02932_),
    .A2(_02934_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08270_ (.A1(_02719_),
    .A2(_02931_),
    .B(_02935_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08271_ (.A1(_02300_),
    .A2(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08272_ (.A1(\as2650.insin[6] ),
    .A2(_02317_),
    .B(_02151_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08273_ (.A1(_02937_),
    .A2(_02938_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08274_ (.A1(_02729_),
    .A2(_02931_),
    .B(_02935_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08275_ (.A1(_02300_),
    .A2(_02939_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08276_ (.A1(\as2650.insin[7] ),
    .A2(_02317_),
    .B(_02151_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08277_ (.A1(_02940_),
    .A2(_02941_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08278_ (.A1(_01272_),
    .A2(_01532_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08279_ (.I(_02162_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08280_ (.A1(_02934_),
    .A2(_02942_),
    .A3(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08281_ (.I(_02944_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08282_ (.I(_02945_),
    .Z(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08283_ (.I(_02945_),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08284_ (.A1(\as2650.ivectors_base[0] ),
    .A2(_02947_),
    .B(_02631_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08285_ (.A1(_01607_),
    .A2(_02946_),
    .B(_02948_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08286_ (.I(_00855_),
    .Z(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08287_ (.A1(\as2650.ivectors_base[1] ),
    .A2(_02947_),
    .B(_02631_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08288_ (.A1(_02949_),
    .A2(_02946_),
    .B(_02950_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08289_ (.I(_00874_),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08290_ (.I(_02630_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08291_ (.A1(\as2650.ivectors_base[2] ),
    .A2(_02947_),
    .B(_02952_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08292_ (.A1(_02951_),
    .A2(_02946_),
    .B(_02953_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08293_ (.I(_01639_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08294_ (.A1(\as2650.ivectors_base[3] ),
    .A2(_02947_),
    .B(_02952_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08295_ (.A1(_02954_),
    .A2(_02946_),
    .B(_02955_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08296_ (.I(_01287_),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08297_ (.I(_02945_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08298_ (.I(_02944_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08299_ (.A1(\as2650.ivectors_base[4] ),
    .A2(_02958_),
    .B(_02952_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08300_ (.A1(_02956_),
    .A2(_02957_),
    .B(_02959_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08301_ (.A1(\as2650.ivectors_base[5] ),
    .A2(_02958_),
    .B(_02952_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08302_ (.A1(_00749_),
    .A2(_02957_),
    .B(_02960_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08303_ (.I(_02630_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08304_ (.A1(\as2650.ivectors_base[6] ),
    .A2(_02958_),
    .B(_02961_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08305_ (.A1(_00772_),
    .A2(_02957_),
    .B(_02962_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08306_ (.A1(\as2650.ivectors_base[7] ),
    .A2(_02958_),
    .B(_02961_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08307_ (.A1(_00796_),
    .A2(_02957_),
    .B(_02963_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08308_ (.I(_02945_),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08309_ (.I(_02944_),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08310_ (.A1(\as2650.ivectors_base[8] ),
    .A2(_02965_),
    .B(_02961_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08311_ (.A1(_00822_),
    .A2(_02964_),
    .B(_02966_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _08312_ (.I(net192),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08313_ (.A1(\as2650.ivectors_base[9] ),
    .A2(_02965_),
    .B(_02961_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08314_ (.A1(_02967_),
    .A2(_02964_),
    .B(_02968_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08315_ (.I(_00879_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08316_ (.I(_01550_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08317_ (.I(_02970_),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08318_ (.A1(\as2650.ivectors_base[10] ),
    .A2(_02965_),
    .B(_02971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08319_ (.A1(_02969_),
    .A2(_02964_),
    .B(_02972_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08320_ (.A1(\as2650.ivectors_base[11] ),
    .A2(_02965_),
    .B(_02971_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08321_ (.A1(_00699_),
    .A2(_02964_),
    .B(_02973_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08322_ (.I(_01150_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08323_ (.A1(_01270_),
    .A2(_01383_),
    .Z(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08324_ (.A1(_02660_),
    .A2(_01258_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08325_ (.I(_02234_),
    .Z(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08326_ (.I(_02977_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08327_ (.I(_02183_),
    .Z(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08328_ (.I(\as2650.stack[0][0] ),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08329_ (.A1(_02847_),
    .A2(_02980_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08330_ (.A1(_02978_),
    .A2(\as2650.stack[1][0] ),
    .B(_02979_),
    .C(_02981_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08331_ (.I(_02196_),
    .Z(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08332_ (.A1(\as2650.stack[3][0] ),
    .A2(_02983_),
    .B1(_02860_),
    .B2(\as2650.stack[2][0] ),
    .C(_02209_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08333_ (.I(\as2650.stack[4][0] ),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08334_ (.A1(_01838_),
    .A2(_02985_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08335_ (.A1(_02978_),
    .A2(\as2650.stack[5][0] ),
    .B(_02979_),
    .C(_02986_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08336_ (.I(_02219_),
    .Z(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08337_ (.A1(\as2650.stack[7][0] ),
    .A2(_02983_),
    .B1(_02860_),
    .B2(\as2650.stack[6][0] ),
    .C(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08338_ (.A1(_02982_),
    .A2(_02984_),
    .B1(_02987_),
    .B2(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08339_ (.I(\as2650.stack[8][0] ),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08340_ (.A1(_02847_),
    .A2(_02991_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08341_ (.A1(_02978_),
    .A2(\as2650.stack[9][0] ),
    .B(_02979_),
    .C(_02992_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08342_ (.A1(\as2650.stack[11][0] ),
    .A2(_02983_),
    .B1(_02202_),
    .B2(\as2650.stack[10][0] ),
    .C(_02209_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08343_ (.I(\as2650.stack[12][0] ),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08344_ (.A1(_01838_),
    .A2(_02995_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08345_ (.A1(_02978_),
    .A2(\as2650.stack[13][0] ),
    .B(_02979_),
    .C(_02996_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08346_ (.A1(\as2650.stack[15][0] ),
    .A2(_02983_),
    .B1(_02860_),
    .B2(\as2650.stack[14][0] ),
    .C(_02988_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08347_ (.A1(_02993_),
    .A2(_02994_),
    .B1(_02997_),
    .B2(_02998_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08348_ (.I0(_02990_),
    .I1(_02999_),
    .S(_02252_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08349_ (.A1(_01397_),
    .A2(_01369_),
    .A3(_03000_),
    .B(_01270_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08350_ (.A1(_02975_),
    .A2(_02976_),
    .A3(_03001_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08351_ (.A1(_02974_),
    .A2(_03002_),
    .B(_02360_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08352_ (.I(_03000_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08353_ (.A1(_01397_),
    .A2(_01369_),
    .A3(_03004_),
    .B(_01270_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08354_ (.A1(_02975_),
    .A2(_02976_),
    .A3(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08355_ (.A1(_02360_),
    .A2(_01151_),
    .A3(_03006_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08356_ (.I(_02833_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08357_ (.A1(_00630_),
    .A2(_03008_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08358_ (.A1(_01653_),
    .A2(_03009_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08359_ (.I(_03010_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08360_ (.A1(_03003_),
    .A2(_03007_),
    .B(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08361_ (.A1(_02705_),
    .A2(_01171_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08362_ (.A1(_00944_),
    .A2(_03013_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08363_ (.I(_03014_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08364_ (.I(_02834_),
    .Z(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08365_ (.A1(_01042_),
    .A2(_02835_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08366_ (.I(_01654_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08367_ (.A1(_03016_),
    .A2(_02362_),
    .B(_03017_),
    .C(_03018_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08368_ (.A1(_03012_),
    .A2(_03015_),
    .A3(_03019_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08369_ (.I(_02789_),
    .Z(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08370_ (.A1(_02360_),
    .A2(_03021_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08371_ (.A1(_02371_),
    .A2(_03014_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08372_ (.I(_03023_),
    .Z(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08373_ (.A1(_03022_),
    .A2(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08374_ (.A1(_02352_),
    .A2(net204),
    .A3(_02796_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08375_ (.A1(net204),
    .A2(_02796_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08376_ (.A1(_02347_),
    .A2(_03027_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08377_ (.A1(_03026_),
    .A2(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08378_ (.I(_02791_),
    .Z(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08379_ (.A1(_03020_),
    .A2(_03025_),
    .B1(_03029_),
    .B2(_03030_),
    .C(_02574_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08380_ (.A1(_03026_),
    .A2(_02808_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08381_ (.I(_02789_),
    .Z(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08382_ (.I(_00944_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08383_ (.A1(_03033_),
    .A2(_02386_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08384_ (.A1(_03032_),
    .A2(_03034_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08385_ (.I(_03008_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08386_ (.A1(_03036_),
    .A2(_03034_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08387_ (.A1(_03016_),
    .A2(_02391_),
    .B(_03037_),
    .C(_01654_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08388_ (.I(_02259_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08389_ (.A1(_01383_),
    .A2(_03039_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08390_ (.I(\as2650.stack[0][1] ),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08391_ (.A1(_02849_),
    .A2(_03041_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08392_ (.A1(_02190_),
    .A2(\as2650.stack[1][1] ),
    .B(_02844_),
    .C(_03042_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08393_ (.I(_02197_),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08394_ (.I(_02861_),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08395_ (.A1(\as2650.stack[3][1] ),
    .A2(_03044_),
    .B1(_03045_),
    .B2(\as2650.stack[2][1] ),
    .C(_02865_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08396_ (.I(_02237_),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08397_ (.I(_02184_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08398_ (.I(\as2650.stack[4][1] ),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08399_ (.A1(_02175_),
    .A2(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08400_ (.A1(_03047_),
    .A2(\as2650.stack[5][1] ),
    .B(_03048_),
    .C(_03050_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08401_ (.A1(\as2650.stack[7][1] ),
    .A2(_02857_),
    .B1(_03045_),
    .B2(\as2650.stack[6][1] ),
    .C(_02221_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08402_ (.A1(_03043_),
    .A2(_03046_),
    .B1(_03051_),
    .B2(_03052_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08403_ (.I(\as2650.stack[8][1] ),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08404_ (.A1(_02175_),
    .A2(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08405_ (.A1(_02190_),
    .A2(\as2650.stack[9][1] ),
    .B(_03048_),
    .C(_03055_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08406_ (.A1(\as2650.stack[11][1] ),
    .A2(_03044_),
    .B1(_03045_),
    .B2(\as2650.stack[10][1] ),
    .C(_02210_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08407_ (.I(\as2650.stack[12][1] ),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08408_ (.A1(_02175_),
    .A2(_03058_),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08409_ (.A1(_03047_),
    .A2(\as2650.stack[13][1] ),
    .B(_03048_),
    .C(_03059_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08410_ (.A1(\as2650.stack[15][1] ),
    .A2(_03044_),
    .B1(_03045_),
    .B2(\as2650.stack[14][1] ),
    .C(_02221_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08411_ (.A1(_03056_),
    .A2(_03057_),
    .B1(_03060_),
    .B2(_03061_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08412_ (.I0(_03053_),
    .I1(_03062_),
    .S(_02253_),
    .Z(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08413_ (.I(_03039_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08414_ (.I(_02430_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08415_ (.A1(_02350_),
    .A2(_01163_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08416_ (.A1(_03065_),
    .A2(_03066_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08417_ (.A1(_02351_),
    .A2(_02430_),
    .A3(_01250_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08418_ (.A1(_01383_),
    .A2(_03067_),
    .A3(_03068_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08419_ (.A1(_02386_),
    .A2(_03040_),
    .B1(_03063_),
    .B2(_03064_),
    .C(_03069_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08420_ (.A1(_01151_),
    .A2(_03070_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08421_ (.A1(_02430_),
    .A2(_02173_),
    .B(_03010_),
    .C(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08422_ (.A1(_03038_),
    .A2(_03072_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08423_ (.A1(_03013_),
    .A2(_03035_),
    .B1(_03073_),
    .B2(_03015_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08424_ (.A1(_02793_),
    .A2(_03031_),
    .B(_03074_),
    .C(_02901_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08425_ (.A1(_03033_),
    .A2(_02413_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08426_ (.A1(_03021_),
    .A2(_03075_),
    .B(_02790_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08427_ (.A1(_02835_),
    .A2(_03075_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08428_ (.A1(_03016_),
    .A2(_02419_),
    .B(_03077_),
    .C(_02606_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08429_ (.I(_02410_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08430_ (.I(_03010_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08431_ (.A1(_01382_),
    .A2(_02260_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08432_ (.I(_03081_),
    .Z(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08433_ (.A1(_02413_),
    .A2(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08434_ (.A1(_03079_),
    .A2(_03067_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08435_ (.I(\as2650.stack[0][2] ),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08436_ (.A1(_02236_),
    .A2(_03085_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08437_ (.A1(_01839_),
    .A2(\as2650.stack[1][2] ),
    .B(_02184_),
    .C(_03086_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08438_ (.I(_02202_),
    .Z(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08439_ (.I(_02209_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08440_ (.A1(\as2650.stack[3][2] ),
    .A2(_02855_),
    .B1(_03088_),
    .B2(\as2650.stack[2][2] ),
    .C(_03089_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08441_ (.I(\as2650.stack[4][2] ),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08442_ (.A1(_02236_),
    .A2(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08443_ (.A1(_02188_),
    .A2(\as2650.stack[5][2] ),
    .B(_02842_),
    .C(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08444_ (.A1(\as2650.stack[7][2] ),
    .A2(_02197_),
    .B1(_03088_),
    .B2(\as2650.stack[6][2] ),
    .C(_02988_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08445_ (.A1(_03087_),
    .A2(_03090_),
    .B1(_03093_),
    .B2(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08446_ (.I(\as2650.stack[8][2] ),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08447_ (.A1(_02236_),
    .A2(_03096_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08448_ (.A1(_02188_),
    .A2(\as2650.stack[9][2] ),
    .B(_02842_),
    .C(_03097_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08449_ (.A1(\as2650.stack[11][2] ),
    .A2(_02855_),
    .B1(_03088_),
    .B2(\as2650.stack[10][2] ),
    .C(_03089_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08450_ (.I(\as2650.stack[12][2] ),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08451_ (.A1(_02847_),
    .A2(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08452_ (.A1(_02188_),
    .A2(\as2650.stack[13][2] ),
    .B(_02842_),
    .C(_03101_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08453_ (.A1(\as2650.stack[15][2] ),
    .A2(_02855_),
    .B1(_03088_),
    .B2(\as2650.stack[14][2] ),
    .C(_02988_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08454_ (.A1(_03098_),
    .A2(_03099_),
    .B1(_03102_),
    .B2(_03103_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08455_ (.I0(_03095_),
    .I1(_03104_),
    .S(_02252_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08456_ (.A1(_01384_),
    .A2(_03084_),
    .B1(_03105_),
    .B2(_02831_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08457_ (.A1(_02974_),
    .A2(_03083_),
    .A3(_03106_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08458_ (.A1(_03079_),
    .A2(_02316_),
    .B(_03080_),
    .C(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08459_ (.A1(_00931_),
    .A2(_02790_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08460_ (.I(_03109_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08461_ (.A1(_03078_),
    .A2(_03108_),
    .B(_03110_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08462_ (.A1(_02806_),
    .A2(_02809_),
    .A3(_02810_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08463_ (.A1(_02811_),
    .A2(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08464_ (.A1(_03076_),
    .A2(_03111_),
    .B1(_03113_),
    .B2(_02372_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08465_ (.A1(_02725_),
    .A2(_03114_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08466_ (.A1(_00632_),
    .A2(_02318_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08467_ (.A1(_02410_),
    .A2(_02429_),
    .A3(_03067_),
    .Z(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08468_ (.A1(_03079_),
    .A2(_03067_),
    .B(_02429_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08469_ (.A1(_03116_),
    .A2(_03117_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08470_ (.I(_01840_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08471_ (.I(\as2650.stack[0][3] ),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08472_ (.A1(_03047_),
    .A2(_03120_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08473_ (.A1(_03119_),
    .A2(\as2650.stack[1][3] ),
    .B(_02186_),
    .C(_03121_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08474_ (.I(_02204_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08475_ (.A1(\as2650.stack[3][3] ),
    .A2(_02199_),
    .B1(_03123_),
    .B2(\as2650.stack[2][3] ),
    .C(_02211_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08476_ (.I(\as2650.stack[4][3] ),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08477_ (.A1(_02238_),
    .A2(_03125_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08478_ (.A1(_03119_),
    .A2(\as2650.stack[5][3] ),
    .B(_02186_),
    .C(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08479_ (.A1(\as2650.stack[7][3] ),
    .A2(_02199_),
    .B1(_03123_),
    .B2(\as2650.stack[6][3] ),
    .C(_02222_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08480_ (.A1(_03122_),
    .A2(_03124_),
    .B1(_03127_),
    .B2(_03128_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08481_ (.I(\as2650.stack[8][3] ),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08482_ (.A1(_03047_),
    .A2(_03130_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08483_ (.A1(_03119_),
    .A2(\as2650.stack[9][3] ),
    .B(_02186_),
    .C(_03131_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08484_ (.I(_02861_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08485_ (.A1(\as2650.stack[11][3] ),
    .A2(_02229_),
    .B1(_03133_),
    .B2(\as2650.stack[10][3] ),
    .C(_02211_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08486_ (.I(_01840_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08487_ (.I(_02185_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08488_ (.I(\as2650.stack[12][3] ),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08489_ (.A1(_02238_),
    .A2(_03137_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08490_ (.A1(_03135_),
    .A2(\as2650.stack[13][3] ),
    .B(_03136_),
    .C(_03138_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08491_ (.A1(\as2650.stack[15][3] ),
    .A2(_02199_),
    .B1(_03123_),
    .B2(\as2650.stack[14][3] ),
    .C(_02243_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08492_ (.A1(_03132_),
    .A2(_03134_),
    .B1(_03139_),
    .B2(_03140_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08493_ (.I0(_03129_),
    .I1(_03141_),
    .S(_02254_),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08494_ (.A1(_01384_),
    .A2(_03118_),
    .B1(_03142_),
    .B2(_02261_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08495_ (.A1(_02433_),
    .A2(_03040_),
    .B(_03143_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08496_ (.A1(_02173_),
    .A2(_03144_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08497_ (.A1(_03011_),
    .A2(_03145_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08498_ (.A1(_01452_),
    .A2(_01398_),
    .A3(_01453_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08499_ (.I(_03147_),
    .Z(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08500_ (.I(_00931_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08501_ (.A1(_03149_),
    .A2(_03148_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08502_ (.A1(_03148_),
    .A2(_02440_),
    .B1(_03150_),
    .B2(_02433_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08503_ (.A1(_03115_),
    .A2(_03146_),
    .B1(_03151_),
    .B2(_01651_),
    .C(_03014_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08504_ (.I(_01457_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08505_ (.I(_03023_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08506_ (.A1(_03153_),
    .A2(_02454_),
    .B(_03154_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08507_ (.A1(_02805_),
    .A2(_02811_),
    .A3(_02814_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08508_ (.A1(_02815_),
    .A2(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08509_ (.I(_02573_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08510_ (.A1(_03152_),
    .A2(_03155_),
    .B1(_03157_),
    .B2(_03030_),
    .C(_03158_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08511_ (.A1(_02803_),
    .A2(_02815_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08512_ (.A1(_02816_),
    .A2(_03159_),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08513_ (.A1(_03021_),
    .A2(_02472_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08514_ (.I(_02451_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08515_ (.I(_03081_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08516_ (.A1(_02453_),
    .A2(_03163_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08517_ (.I(_01382_),
    .Z(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08518_ (.A1(_03162_),
    .A2(_03116_),
    .Z(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08519_ (.I(_02237_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08520_ (.I(\as2650.stack[0][4] ),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08521_ (.A1(_03167_),
    .A2(_03168_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08522_ (.A1(_03135_),
    .A2(\as2650.stack[1][4] ),
    .B(_03136_),
    .C(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08523_ (.A1(\as2650.stack[3][4] ),
    .A2(_02857_),
    .B1(_02862_),
    .B2(\as2650.stack[2][4] ),
    .C(_02865_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08524_ (.I(\as2650.stack[4][4] ),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08525_ (.A1(_03167_),
    .A2(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08526_ (.A1(_03135_),
    .A2(\as2650.stack[5][4] ),
    .B(_02844_),
    .C(_03173_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08527_ (.A1(\as2650.stack[7][4] ),
    .A2(_02229_),
    .B1(_03133_),
    .B2(\as2650.stack[6][4] ),
    .C(_02243_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08528_ (.A1(_03170_),
    .A2(_03171_),
    .B1(_03174_),
    .B2(_03175_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08529_ (.I(\as2650.stack[8][4] ),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08530_ (.A1(_03167_),
    .A2(_03177_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08531_ (.A1(_03135_),
    .A2(\as2650.stack[9][4] ),
    .B(_03136_),
    .C(_03178_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08532_ (.A1(\as2650.stack[11][4] ),
    .A2(_02857_),
    .B1(_02862_),
    .B2(\as2650.stack[10][4] ),
    .C(_02865_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08533_ (.I(\as2650.stack[12][4] ),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08534_ (.A1(_02849_),
    .A2(_03181_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08535_ (.A1(_01841_),
    .A2(\as2650.stack[13][4] ),
    .B(_02844_),
    .C(_03182_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08536_ (.A1(\as2650.stack[15][4] ),
    .A2(_02229_),
    .B1(_03133_),
    .B2(\as2650.stack[14][4] ),
    .C(_02243_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08537_ (.A1(_03179_),
    .A2(_03180_),
    .B1(_03183_),
    .B2(_03184_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08538_ (.I0(_03176_),
    .I1(_03185_),
    .S(_02253_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08539_ (.I(_02260_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08540_ (.A1(_03165_),
    .A2(_03166_),
    .B1(_03186_),
    .B2(_03187_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08541_ (.A1(_03164_),
    .A2(_03188_),
    .B(_02171_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08542_ (.A1(_03162_),
    .A2(_02334_),
    .B(_03189_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08543_ (.A1(_00944_),
    .A2(_03008_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08544_ (.I(_03191_),
    .Z(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08545_ (.A1(_03036_),
    .A2(_02459_),
    .B1(_03192_),
    .B2(_02453_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08546_ (.I(_02266_),
    .Z(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08547_ (.A1(_03080_),
    .A2(_03190_),
    .B1(_03193_),
    .B2(_03194_),
    .C(_03110_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08548_ (.A1(_03024_),
    .A2(_03161_),
    .B(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08549_ (.A1(_02793_),
    .A2(_03160_),
    .B(_03196_),
    .C(_02901_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08550_ (.A1(_02802_),
    .A2(_02817_),
    .A3(_02819_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08551_ (.A1(_02820_),
    .A2(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08552_ (.A1(_03032_),
    .A2(_02494_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08553_ (.I(_02468_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08554_ (.A1(_02470_),
    .A2(_03163_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08555_ (.A1(_02451_),
    .A2(_03200_),
    .A3(_03116_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08556_ (.A1(_03162_),
    .A2(_03116_),
    .B(_03200_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08557_ (.A1(_03202_),
    .A2(_03203_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08558_ (.I(\as2650.stack[0][5] ),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08559_ (.A1(_02848_),
    .A2(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08560_ (.A1(_02189_),
    .A2(\as2650.stack[1][5] ),
    .B(_02843_),
    .C(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08561_ (.A1(\as2650.stack[3][5] ),
    .A2(_02856_),
    .B1(_02203_),
    .B2(\as2650.stack[2][5] ),
    .C(_03089_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08562_ (.I(\as2650.stack[4][5] ),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08563_ (.A1(_02848_),
    .A2(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08564_ (.A1(_02189_),
    .A2(\as2650.stack[5][5] ),
    .B(_02843_),
    .C(_03210_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08565_ (.A1(\as2650.stack[7][5] ),
    .A2(_02856_),
    .B1(_02861_),
    .B2(\as2650.stack[6][5] ),
    .C(_02220_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08566_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03211_),
    .B2(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08567_ (.I(\as2650.stack[8][5] ),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08568_ (.A1(_02848_),
    .A2(_03214_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08569_ (.A1(_02189_),
    .A2(\as2650.stack[9][5] ),
    .B(_02843_),
    .C(_03215_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08570_ (.A1(\as2650.stack[11][5] ),
    .A2(_02197_),
    .B1(_02203_),
    .B2(\as2650.stack[10][5] ),
    .C(_03089_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08571_ (.I(\as2650.stack[12][5] ),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08572_ (.A1(_01839_),
    .A2(_03218_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08573_ (.A1(_02237_),
    .A2(\as2650.stack[13][5] ),
    .B(_02184_),
    .C(_03219_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08574_ (.A1(\as2650.stack[15][5] ),
    .A2(_02856_),
    .B1(_02203_),
    .B2(\as2650.stack[14][5] ),
    .C(_02220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08575_ (.A1(_03216_),
    .A2(_03217_),
    .B1(_03220_),
    .B2(_03221_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08576_ (.I0(_03213_),
    .I1(_03222_),
    .S(_02253_),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08577_ (.A1(_03165_),
    .A2(_03204_),
    .B1(_03223_),
    .B2(_03187_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08578_ (.A1(_03201_),
    .A2(_03224_),
    .B(_02298_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08579_ (.A1(_03200_),
    .A2(_02334_),
    .B(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08580_ (.I(_03147_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08581_ (.A1(_03227_),
    .A2(_02477_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08582_ (.A1(_02470_),
    .A2(_03192_),
    .B(_03228_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08583_ (.A1(_03080_),
    .A2(_03226_),
    .B1(_03229_),
    .B2(_03194_),
    .C(_03110_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08584_ (.A1(_03024_),
    .A2(_03199_),
    .B(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08585_ (.A1(_02792_),
    .A2(_03198_),
    .B(_03231_),
    .C(_02901_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08586_ (.I(_02510_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08587_ (.I(_02298_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08588_ (.I(_02492_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08589_ (.A1(_03234_),
    .A2(_03082_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08590_ (.I(_01382_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08591_ (.A1(_03232_),
    .A2(_03202_),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08592_ (.I(\as2650.stack[0][6] ),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08593_ (.A1(_02235_),
    .A2(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08594_ (.A1(_02977_),
    .A2(\as2650.stack[1][6] ),
    .B(_02183_),
    .C(_03239_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08595_ (.I(_02201_),
    .Z(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08596_ (.A1(\as2650.stack[3][6] ),
    .A2(_02195_),
    .B1(_03241_),
    .B2(\as2650.stack[2][6] ),
    .C(_02208_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08597_ (.I(\as2650.stack[4][6] ),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08598_ (.A1(_01837_),
    .A2(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08599_ (.A1(_02977_),
    .A2(\as2650.stack[5][6] ),
    .B(_02182_),
    .C(_03244_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08600_ (.A1(\as2650.stack[7][6] ),
    .A2(_02196_),
    .B1(_03241_),
    .B2(\as2650.stack[6][6] ),
    .C(_02219_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08601_ (.A1(_03240_),
    .A2(_03242_),
    .B1(_03245_),
    .B2(_03246_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08602_ (.I(\as2650.stack[8][6] ),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08603_ (.A1(_01837_),
    .A2(_03248_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08604_ (.A1(_02977_),
    .A2(\as2650.stack[9][6] ),
    .B(_02182_),
    .C(_03249_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08605_ (.A1(\as2650.stack[11][6] ),
    .A2(_02195_),
    .B1(_03241_),
    .B2(\as2650.stack[10][6] ),
    .C(_02208_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08606_ (.I(\as2650.stack[12][6] ),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08607_ (.A1(_01837_),
    .A2(_03252_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08608_ (.A1(_02235_),
    .A2(\as2650.stack[13][6] ),
    .B(_02182_),
    .C(_03253_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08609_ (.A1(\as2650.stack[15][6] ),
    .A2(_02195_),
    .B1(_03241_),
    .B2(\as2650.stack[14][6] ),
    .C(_02219_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08610_ (.A1(_03250_),
    .A2(_03251_),
    .B1(_03254_),
    .B2(_03255_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08611_ (.I0(_03247_),
    .I1(_03256_),
    .S(_02252_),
    .Z(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08612_ (.A1(_03236_),
    .A2(_03237_),
    .B1(_03257_),
    .B2(_03187_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08613_ (.A1(_03235_),
    .A2(_03258_),
    .B(_02171_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08614_ (.A1(_03232_),
    .A2(_03233_),
    .B(_03259_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08615_ (.A1(_02357_),
    .A2(_02497_),
    .B(_02500_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08616_ (.A1(_03234_),
    .A2(_03192_),
    .B1(_03261_),
    .B2(_02835_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08617_ (.A1(_03011_),
    .A2(_03260_),
    .B1(_03262_),
    .B2(_03018_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08618_ (.A1(_03015_),
    .A2(_03263_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08619_ (.A1(_03153_),
    .A2(_03234_),
    .B(_03154_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08620_ (.A1(_02800_),
    .A2(_02820_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08621_ (.A1(_02821_),
    .A2(_03266_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08622_ (.A1(_03264_),
    .A2(_03265_),
    .B1(_03267_),
    .B2(_03030_),
    .C(_03158_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08623_ (.A1(_02799_),
    .A2(_02822_),
    .A3(_02824_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08624_ (.A1(_02825_),
    .A2(_03268_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08625_ (.A1(_03032_),
    .A2(_02513_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08626_ (.I(\as2650.PC[7] ),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08627_ (.A1(_02514_),
    .A2(_03163_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08628_ (.A1(_02510_),
    .A2(_03271_),
    .A3(_03202_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08629_ (.A1(_03232_),
    .A2(_03202_),
    .B(_03271_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08630_ (.A1(_03273_),
    .A2(_03274_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08631_ (.I(_02181_),
    .Z(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08632_ (.I(\as2650.stack[0][7] ),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08633_ (.A1(_01836_),
    .A2(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08634_ (.A1(_02234_),
    .A2(\as2650.stack[1][7] ),
    .B(_03276_),
    .C(_03278_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08635_ (.I(_02179_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08636_ (.A1(\as2650.stack[3][7] ),
    .A2(_03280_),
    .B1(_02180_),
    .B2(\as2650.stack[2][7] ),
    .C(_02208_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08637_ (.I(\as2650.stack[4][7] ),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08638_ (.A1(_02233_),
    .A2(_03282_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08639_ (.A1(_01836_),
    .A2(\as2650.stack[5][7] ),
    .B(_03276_),
    .C(_03283_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08640_ (.A1(\as2650.stack[7][7] ),
    .A2(_03280_),
    .B1(_02201_),
    .B2(\as2650.stack[6][7] ),
    .C(_02218_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08641_ (.A1(_03279_),
    .A2(_03281_),
    .B1(_03284_),
    .B2(_03285_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08642_ (.I(\as2650.stack[8][7] ),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08643_ (.A1(_02233_),
    .A2(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08644_ (.A1(_02234_),
    .A2(\as2650.stack[9][7] ),
    .B(_03276_),
    .C(_03288_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08645_ (.A1(\as2650.stack[11][7] ),
    .A2(_03280_),
    .B1(_02180_),
    .B2(\as2650.stack[10][7] ),
    .C(_02207_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08646_ (.I(\as2650.stack[12][7] ),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08647_ (.A1(_02233_),
    .A2(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08648_ (.A1(_01836_),
    .A2(\as2650.stack[13][7] ),
    .B(_03276_),
    .C(_03292_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08649_ (.A1(\as2650.stack[15][7] ),
    .A2(_03280_),
    .B1(_02201_),
    .B2(\as2650.stack[14][7] ),
    .C(_02218_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08650_ (.A1(_03289_),
    .A2(_03290_),
    .B1(_03293_),
    .B2(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08651_ (.I0(_03286_),
    .I1(_03295_),
    .S(_02251_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08652_ (.A1(_03165_),
    .A2(_03275_),
    .B1(_03296_),
    .B2(_03039_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08653_ (.A1(_03272_),
    .A2(_03297_),
    .B(_02298_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08654_ (.A1(_03271_),
    .A2(_02334_),
    .B(_03298_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08655_ (.A1(_03036_),
    .A2(_02518_),
    .B1(_03192_),
    .B2(_02514_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08656_ (.A1(_03080_),
    .A2(_03299_),
    .B1(_03300_),
    .B2(_03194_),
    .C(_03110_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08657_ (.A1(_03154_),
    .A2(_03270_),
    .B(_03301_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08658_ (.I(_01080_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08659_ (.A1(_02792_),
    .A2(_03269_),
    .B(_03302_),
    .C(_03303_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08660_ (.I(_02547_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08661_ (.A1(_02355_),
    .A2(_02533_),
    .B(_02499_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08662_ (.A1(_03304_),
    .A2(_03191_),
    .B1(_03305_),
    .B2(_03008_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08663_ (.I(_02528_),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08664_ (.A1(_03304_),
    .A2(_03163_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08665_ (.A1(_03307_),
    .A2(_03273_),
    .Z(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08666_ (.I(_02238_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08667_ (.I(_02185_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08668_ (.I(_01840_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08669_ (.I(\as2650.stack[0][8] ),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08670_ (.A1(_03312_),
    .A2(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08671_ (.A1(_03310_),
    .A2(\as2650.stack[1][8] ),
    .B(_03311_),
    .C(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08672_ (.I(_02210_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08673_ (.A1(\as2650.stack[3][8] ),
    .A2(_02914_),
    .B1(_02205_),
    .B2(\as2650.stack[2][8] ),
    .C(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08674_ (.I(_02185_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08675_ (.I(\as2650.stack[4][8] ),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08676_ (.A1(_03312_),
    .A2(_03319_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08677_ (.A1(_03310_),
    .A2(\as2650.stack[5][8] ),
    .B(_03318_),
    .C(_03320_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08678_ (.I(_02198_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08679_ (.I(_02204_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08680_ (.A1(\as2650.stack[7][8] ),
    .A2(_03322_),
    .B1(_03323_),
    .B2(\as2650.stack[6][8] ),
    .C(_02222_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08681_ (.A1(_03315_),
    .A2(_03317_),
    .B1(_03321_),
    .B2(_03324_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08682_ (.I(\as2650.stack[8][8] ),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08683_ (.A1(_03312_),
    .A2(_03326_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08684_ (.A1(_03310_),
    .A2(\as2650.stack[9][8] ),
    .B(_03318_),
    .C(_03327_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08685_ (.A1(\as2650.stack[11][8] ),
    .A2(_02914_),
    .B1(_02205_),
    .B2(\as2650.stack[10][8] ),
    .C(_02211_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08686_ (.I(_03167_),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08687_ (.I(\as2650.stack[12][8] ),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08688_ (.A1(_03119_),
    .A2(_03331_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08689_ (.A1(_03330_),
    .A2(\as2650.stack[13][8] ),
    .B(_03318_),
    .C(_03332_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08690_ (.A1(\as2650.stack[15][8] ),
    .A2(_02914_),
    .B1(_03323_),
    .B2(\as2650.stack[14][8] ),
    .C(_02222_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08691_ (.A1(_03328_),
    .A2(_03329_),
    .B1(_03333_),
    .B2(_03334_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08692_ (.I0(_03325_),
    .I1(_03335_),
    .S(_02254_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08693_ (.A1(_03165_),
    .A2(_03309_),
    .B1(_03336_),
    .B2(_03039_),
    .C(_01647_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08694_ (.A1(_02737_),
    .A2(_03306_),
    .B1(_03308_),
    .B2(_03337_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08695_ (.A1(_03307_),
    .A2(_02974_),
    .B1(_03338_),
    .B2(_01488_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08696_ (.A1(_03011_),
    .A2(_03306_),
    .B(_03339_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08697_ (.A1(_03015_),
    .A2(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08698_ (.A1(_03153_),
    .A2(_03304_),
    .B(_03154_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08699_ (.A1(_02797_),
    .A2(_02825_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08700_ (.A1(_00899_),
    .A2(_03343_),
    .Z(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08701_ (.A1(_03341_),
    .A2(_03342_),
    .B1(_03344_),
    .B2(_03030_),
    .C(_03158_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08702_ (.I(_02543_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08703_ (.A1(_02737_),
    .A2(_03009_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08704_ (.I(_02545_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08705_ (.A1(_03347_),
    .A2(_03081_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08706_ (.A1(_03307_),
    .A2(_03273_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08707_ (.A1(_03345_),
    .A2(_03349_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08708_ (.I(_03048_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08709_ (.I(\as2650.stack[0][9] ),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08710_ (.A1(_02176_),
    .A2(_03352_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08711_ (.A1(_02239_),
    .A2(\as2650.stack[1][9] ),
    .B(_03351_),
    .C(_03353_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08712_ (.A1(\as2650.stack[3][9] ),
    .A2(_03322_),
    .B1(_03323_),
    .B2(\as2650.stack[2][9] ),
    .C(_03316_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08713_ (.I(\as2650.stack[4][9] ),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08714_ (.A1(_02176_),
    .A2(_03356_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08715_ (.A1(_02239_),
    .A2(\as2650.stack[5][9] ),
    .B(_03311_),
    .C(_03357_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08716_ (.I(_03044_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08717_ (.I(_02204_),
    .Z(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08718_ (.I(_02221_),
    .Z(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08719_ (.A1(\as2650.stack[7][9] ),
    .A2(_03359_),
    .B1(_03360_),
    .B2(\as2650.stack[6][9] ),
    .C(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08720_ (.A1(_03354_),
    .A2(_03355_),
    .B1(_03358_),
    .B2(_03362_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08721_ (.I(\as2650.stack[8][9] ),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08722_ (.A1(_02176_),
    .A2(_03364_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08723_ (.A1(_02239_),
    .A2(\as2650.stack[9][9] ),
    .B(_03311_),
    .C(_03365_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08724_ (.A1(\as2650.stack[11][9] ),
    .A2(_03322_),
    .B1(_03323_),
    .B2(\as2650.stack[10][9] ),
    .C(_03316_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08725_ (.I(\as2650.stack[12][9] ),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08726_ (.A1(_03312_),
    .A2(_03368_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08727_ (.A1(_03310_),
    .A2(\as2650.stack[13][9] ),
    .B(_03311_),
    .C(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08728_ (.A1(\as2650.stack[15][9] ),
    .A2(_03322_),
    .B1(_03360_),
    .B2(\as2650.stack[14][9] ),
    .C(_03361_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08729_ (.A1(_03366_),
    .A2(_03367_),
    .B1(_03370_),
    .B2(_03371_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08730_ (.I0(_03363_),
    .I1(_03372_),
    .S(_02254_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08731_ (.A1(_03236_),
    .A2(_03350_),
    .B1(_03373_),
    .B2(_03187_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08732_ (.A1(_02315_),
    .A2(_03348_),
    .A3(_03374_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08733_ (.A1(_01205_),
    .A2(_03345_),
    .B(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08734_ (.A1(_01376_),
    .A2(_02834_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08735_ (.A1(_00931_),
    .A2(_03347_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08736_ (.A1(_03227_),
    .A2(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08737_ (.A1(_02551_),
    .A2(_03377_),
    .B(_03379_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08738_ (.A1(_03346_),
    .A2(_03376_),
    .B1(_03380_),
    .B2(_03194_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08739_ (.A1(_03345_),
    .A2(_02422_),
    .B(_03014_),
    .C(_03381_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08740_ (.A1(_03153_),
    .A2(_03347_),
    .B(_03023_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08741_ (.A1(_02749_),
    .A2(_02826_),
    .Z(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08742_ (.A1(_03382_),
    .A2(_03383_),
    .B1(_03384_),
    .B2(_02793_),
    .C(_03158_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08743_ (.A1(_02541_),
    .A2(_02826_),
    .B(_02570_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08744_ (.A1(_03149_),
    .A2(_02562_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08745_ (.A1(_03032_),
    .A2(_03386_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08746_ (.A1(_03021_),
    .A2(_02827_),
    .A3(_03385_),
    .B(_03387_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08747_ (.A1(_02568_),
    .A2(_03377_),
    .B1(_03386_),
    .B2(_03036_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08748_ (.A1(_01650_),
    .A2(_03389_),
    .Z(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08749_ (.A1(_02528_),
    .A2(_02543_),
    .A3(_03273_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08750_ (.A1(_02577_),
    .A2(_03391_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08751_ (.I(\as2650.stack[0][10] ),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08752_ (.A1(_02850_),
    .A2(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08753_ (.A1(_02885_),
    .A2(\as2650.stack[1][10] ),
    .B(_02845_),
    .C(_03394_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08754_ (.A1(\as2650.stack[3][10] ),
    .A2(_03359_),
    .B1(_03360_),
    .B2(\as2650.stack[2][10] ),
    .C(_02866_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08755_ (.I(\as2650.stack[4][10] ),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08756_ (.A1(_02917_),
    .A2(_03397_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08757_ (.A1(_02885_),
    .A2(\as2650.stack[5][10] ),
    .B(_03351_),
    .C(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08758_ (.A1(\as2650.stack[7][10] ),
    .A2(_02858_),
    .B1(_02863_),
    .B2(\as2650.stack[6][10] ),
    .C(_03361_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08759_ (.A1(_03395_),
    .A2(_03396_),
    .B1(_03399_),
    .B2(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08760_ (.I(\as2650.stack[8][10] ),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08761_ (.A1(_02917_),
    .A2(_03402_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08762_ (.A1(_02885_),
    .A2(\as2650.stack[9][10] ),
    .B(_03351_),
    .C(_03403_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08763_ (.A1(\as2650.stack[11][10] ),
    .A2(_03359_),
    .B1(_03360_),
    .B2(\as2650.stack[10][10] ),
    .C(_03316_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08764_ (.I(\as2650.stack[12][10] ),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08765_ (.A1(_02917_),
    .A2(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08766_ (.A1(_02191_),
    .A2(\as2650.stack[13][10] ),
    .B(_03351_),
    .C(_03407_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08767_ (.A1(\as2650.stack[15][10] ),
    .A2(_03359_),
    .B1(_02863_),
    .B2(\as2650.stack[14][10] ),
    .C(_03361_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08768_ (.A1(_03404_),
    .A2(_03405_),
    .B1(_03408_),
    .B2(_03409_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08769_ (.I0(_03401_),
    .I1(_03410_),
    .S(_02255_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08770_ (.A1(_03236_),
    .A2(_03392_),
    .B1(_03411_),
    .B2(_02261_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08771_ (.A1(_02562_),
    .A2(_03040_),
    .B(_03412_),
    .C(_02315_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08772_ (.A1(_02558_),
    .A2(_02316_),
    .B(_03010_),
    .C(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08773_ (.A1(_03390_),
    .A2(_03414_),
    .B(_03023_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08774_ (.A1(_03013_),
    .A2(_03388_),
    .B(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08775_ (.A1(_02725_),
    .A2(_03416_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08776_ (.I(_02579_),
    .Z(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08777_ (.A1(_03149_),
    .A2(_01457_),
    .A3(_02790_),
    .A4(_03417_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08778_ (.I(_02576_),
    .Z(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08779_ (.A1(_02577_),
    .A2(_03391_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08780_ (.A1(_02576_),
    .A2(_03420_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08781_ (.A1(_03419_),
    .A2(_03420_),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08782_ (.A1(_01384_),
    .A2(_03421_),
    .A3(_03422_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08783_ (.I(_03136_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08784_ (.I(\as2650.stack[0][11] ),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08785_ (.A1(_03330_),
    .A2(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08786_ (.A1(_02232_),
    .A2(\as2650.stack[1][11] ),
    .B(_03424_),
    .C(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08787_ (.I(_02862_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08788_ (.A1(\as2650.stack[3][11] ),
    .A2(_02230_),
    .B1(_03428_),
    .B2(\as2650.stack[2][11] ),
    .C(_02866_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08789_ (.I(\as2650.stack[4][11] ),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08790_ (.A1(_03330_),
    .A2(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08791_ (.A1(_01842_),
    .A2(\as2650.stack[5][11] ),
    .B(_03424_),
    .C(_03431_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08792_ (.A1(\as2650.stack[7][11] ),
    .A2(_02230_),
    .B1(_03428_),
    .B2(\as2650.stack[6][11] ),
    .C(_02244_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08793_ (.A1(_03427_),
    .A2(_03429_),
    .B1(_03432_),
    .B2(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08794_ (.I(\as2650.stack[8][11] ),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08795_ (.A1(_03330_),
    .A2(_03435_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08796_ (.A1(_02232_),
    .A2(\as2650.stack[9][11] ),
    .B(_03424_),
    .C(_03436_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08797_ (.A1(\as2650.stack[11][11] ),
    .A2(_02858_),
    .B1(_03428_),
    .B2(\as2650.stack[10][11] ),
    .C(_02866_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08798_ (.I(\as2650.stack[12][11] ),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08799_ (.A1(_02850_),
    .A2(_03439_),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08800_ (.A1(_01842_),
    .A2(\as2650.stack[13][11] ),
    .B(_02845_),
    .C(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08801_ (.A1(\as2650.stack[15][11] ),
    .A2(_02230_),
    .B1(_03428_),
    .B2(\as2650.stack[14][11] ),
    .C(_02244_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08802_ (.A1(_03437_),
    .A2(_03438_),
    .B1(_03441_),
    .B2(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08803_ (.I0(_03434_),
    .I1(_03443_),
    .S(_02255_),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08804_ (.A1(_03417_),
    .A2(_03082_),
    .B1(_03444_),
    .B2(_02831_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08805_ (.A1(_01151_),
    .A2(_03423_),
    .A3(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08806_ (.A1(_01206_),
    .A2(_03419_),
    .B(_03446_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08807_ (.A1(_02388_),
    .A2(_03227_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08808_ (.A1(_03149_),
    .A2(_03417_),
    .B(_02834_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08809_ (.A1(_02583_),
    .A2(_03448_),
    .B(_03449_),
    .C(_01654_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08810_ (.A1(_03419_),
    .A2(_01447_),
    .B(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08811_ (.A1(_03346_),
    .A2(_03447_),
    .B(_03451_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08812_ (.A1(\as2650.instruction_args_latch[11] ),
    .A2(_02827_),
    .Z(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08813_ (.A1(_03024_),
    .A2(_03452_),
    .B1(_03453_),
    .B2(_02372_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08814_ (.A1(_02376_),
    .A2(_03418_),
    .A3(_03454_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08815_ (.A1(_02585_),
    .A2(_02827_),
    .B(_02600_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08816_ (.A1(_02897_),
    .A2(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08817_ (.I(_03318_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08818_ (.I(\as2650.stack[0][12] ),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08819_ (.A1(_01842_),
    .A2(_03458_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08820_ (.A1(_02918_),
    .A2(\as2650.stack[1][12] ),
    .B(_03457_),
    .C(_03459_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08821_ (.I(_02205_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08822_ (.A1(\as2650.stack[3][12] ),
    .A2(_02915_),
    .B1(_03461_),
    .B2(\as2650.stack[2][12] ),
    .C(_02212_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08823_ (.I(\as2650.stack[4][12] ),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08824_ (.A1(_02869_),
    .A2(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08825_ (.A1(_02918_),
    .A2(\as2650.stack[5][12] ),
    .B(_03457_),
    .C(_03464_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08826_ (.A1(\as2650.stack[7][12] ),
    .A2(_02915_),
    .B1(_03461_),
    .B2(\as2650.stack[6][12] ),
    .C(_02223_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08827_ (.A1(_03460_),
    .A2(_03462_),
    .B1(_03465_),
    .B2(_03466_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08828_ (.I(\as2650.stack[8][12] ),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08829_ (.A1(_02869_),
    .A2(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08830_ (.A1(_02918_),
    .A2(\as2650.stack[9][12] ),
    .B(_03457_),
    .C(_03469_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08831_ (.A1(\as2650.stack[11][12] ),
    .A2(_02200_),
    .B1(_03461_),
    .B2(\as2650.stack[10][12] ),
    .C(_02212_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08832_ (.I(\as2650.stack[12][12] ),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08833_ (.A1(_02869_),
    .A2(_03472_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08834_ (.A1(_02177_),
    .A2(\as2650.stack[13][12] ),
    .B(_03457_),
    .C(_03473_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08835_ (.A1(\as2650.stack[15][12] ),
    .A2(_02915_),
    .B1(_03461_),
    .B2(\as2650.stack[14][12] ),
    .C(_02223_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08836_ (.A1(_03470_),
    .A2(_03471_),
    .B1(_03474_),
    .B2(_03475_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08837_ (.I0(_03467_),
    .I1(_03476_),
    .S(_02892_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08838_ (.A1(_02596_),
    .A2(_03421_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08839_ (.A1(_03236_),
    .A2(_03478_),
    .Z(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08840_ (.A1(_02598_),
    .A2(_03082_),
    .B1(_03477_),
    .B2(_02831_),
    .C(_03479_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08841_ (.A1(_02596_),
    .A2(_02171_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08842_ (.A1(_02299_),
    .A2(_03480_),
    .B(_03481_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08843_ (.A1(_03033_),
    .A2(_03148_),
    .B1(_03109_),
    .B2(_02606_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08844_ (.A1(_03482_),
    .A2(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08845_ (.A1(_03033_),
    .A2(_02598_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08846_ (.A1(_02789_),
    .A2(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08847_ (.A1(_02599_),
    .A2(_03109_),
    .A3(_03448_),
    .B1(_03485_),
    .B2(_03148_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08848_ (.A1(_03013_),
    .A2(_03486_),
    .B1(_03487_),
    .B2(_03018_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08849_ (.A1(_03484_),
    .A2(_03488_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08850_ (.A1(_02840_),
    .A2(_03456_),
    .B(_03489_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08851_ (.A1(_02725_),
    .A2(_03490_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08852_ (.I(_02696_),
    .Z(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08853_ (.A1(_00938_),
    .A2(_01178_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08854_ (.I(_03492_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08855_ (.A1(_01236_),
    .A2(_01211_),
    .A3(_01260_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08856_ (.A1(_00589_),
    .A2(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _08857_ (.A1(_02257_),
    .A2(_01219_),
    .B(_01255_),
    .C(_03495_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _08858_ (.A1(_01147_),
    .A2(_01433_),
    .A3(_03496_),
    .Z(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08859_ (.I(_03497_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08860_ (.I(_01427_),
    .Z(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08861_ (.I(_01101_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08862_ (.A1(_01300_),
    .A2(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08863_ (.A1(_03500_),
    .A2(_02727_),
    .B(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08864_ (.A1(_01009_),
    .A2(_03500_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08865_ (.A1(_03500_),
    .A2(_01641_),
    .B(_03503_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08866_ (.A1(_03502_),
    .A2(_03504_),
    .Z(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08867_ (.A1(_03502_),
    .A2(_03504_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08868_ (.A1(_03505_),
    .A2(_03506_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08869_ (.I(_01098_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08870_ (.I(_03508_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08871_ (.I(_03509_),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08872_ (.A1(_01312_),
    .A2(_03510_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08873_ (.A1(_01102_),
    .A2(_02490_),
    .B(_03511_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08874_ (.A1(_01013_),
    .A2(_03510_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08875_ (.A1(_03510_),
    .A2(_01631_),
    .B(_03513_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08876_ (.I(_03514_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08877_ (.A1(_03512_),
    .A2(_03515_),
    .Z(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08878_ (.A1(_01092_),
    .A2(_01097_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08879_ (.I(_03517_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08880_ (.I(_03518_),
    .Z(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08881_ (.A1(_03518_),
    .A2(_01134_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08882_ (.A1(_01616_),
    .A2(_03519_),
    .B(_03520_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08883_ (.A1(_01018_),
    .A2(_03510_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08884_ (.A1(_01102_),
    .A2(_01620_),
    .B(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08885_ (.A1(_03521_),
    .A2(_03523_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08886_ (.A1(_03521_),
    .A2(_03523_),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _08887_ (.A1(_03524_),
    .A2(_03525_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08888_ (.A1(_01020_),
    .A2(_01101_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08889_ (.A1(_01101_),
    .A2(_01609_),
    .B(_03527_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08890_ (.I(_03528_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08891_ (.A1(_01329_),
    .A2(_03509_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08892_ (.A1(_03509_),
    .A2(_02447_),
    .B(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08893_ (.I(_03531_),
    .Z(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08894_ (.A1(_03529_),
    .A2(_03532_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08895_ (.I0(_02345_),
    .I1(_01292_),
    .S(_01099_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08896_ (.I(_03517_),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08897_ (.A1(_01466_),
    .A2(_03535_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08898_ (.A1(_01563_),
    .A2(_01304_),
    .B(_03508_),
    .C(_01567_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08899_ (.A1(_03534_),
    .A2(_03536_),
    .A3(_03537_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08900_ (.I(_00726_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08901_ (.A1(_03539_),
    .A2(_03509_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08902_ (.A1(_01628_),
    .A2(_01467_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08903_ (.A1(_01628_),
    .A2(_01359_),
    .B(_03535_),
    .C(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08904_ (.I0(_01086_),
    .I1(_01304_),
    .S(_03508_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08905_ (.A1(_03540_),
    .A2(_03542_),
    .B(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08906_ (.A1(_01517_),
    .A2(\as2650.debug_psl[3] ),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08907_ (.A1(_03538_),
    .A2(_03544_),
    .B(_03545_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08908_ (.A1(_03534_),
    .A2(_03540_),
    .A3(_03542_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08909_ (.A1(_02380_),
    .A2(_03517_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08910_ (.A1(_00760_),
    .A2(_03508_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08911_ (.A1(_03548_),
    .A2(_03549_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(_01474_),
    .A2(_01099_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08913_ (.A1(_01099_),
    .A2(_01579_),
    .B(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08914_ (.I(_03552_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08915_ (.A1(_03550_),
    .A2(_03553_),
    .Z(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08916_ (.A1(_03546_),
    .A2(_03547_),
    .B(_03554_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08917_ (.A1(_03548_),
    .A2(_03549_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(_03556_),
    .A2(_03553_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08919_ (.I(_03557_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08920_ (.A1(_02320_),
    .A2(_03535_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08921_ (.A1(_01338_),
    .A2(_03518_),
    .B(_03559_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08922_ (.A1(_01479_),
    .A2(_01100_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08923_ (.A1(_01100_),
    .A2(_01588_),
    .B(_03561_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08924_ (.A1(_03560_),
    .A2(_03562_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08925_ (.A1(_03560_),
    .A2(_03562_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08926_ (.A1(_03563_),
    .A2(_03564_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08927_ (.A1(_03555_),
    .A2(_03558_),
    .B(_03565_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _08928_ (.A1(_01339_),
    .A2(_03519_),
    .B(_03559_),
    .C(_03562_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08929_ (.A1(_01091_),
    .A2(_03535_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08930_ (.A1(_01284_),
    .A2(_03518_),
    .B(_03568_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08931_ (.A1(_03517_),
    .A2(_01597_),
    .Z(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08932_ (.A1(_00794_),
    .A2(_01100_),
    .B(_03570_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08933_ (.A1(_03569_),
    .A2(_03571_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08934_ (.I(_03572_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08935_ (.A1(_03566_),
    .A2(_03567_),
    .B(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08936_ (.I(_00794_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08937_ (.I(_03569_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08938_ (.A1(_03575_),
    .A2(_01227_),
    .B(_03576_),
    .C(_03570_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08939_ (.A1(_03529_),
    .A2(_03532_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08940_ (.A1(_03533_),
    .A2(_03574_),
    .A3(_03577_),
    .B(_03578_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08941_ (.I(_03521_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08942_ (.A1(_03580_),
    .A2(_03523_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08943_ (.A1(_03526_),
    .A2(_03579_),
    .B(_03581_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08944_ (.I(_03512_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08945_ (.A1(_03583_),
    .A2(_03515_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08946_ (.A1(_03516_),
    .A2(_03582_),
    .B(_03584_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08947_ (.A1(_02156_),
    .A2(_02727_),
    .B(_03501_),
    .C(_03504_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08948_ (.A1(_03507_),
    .A2(_03585_),
    .B(_03586_),
    .C(_01421_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08949_ (.A1(_03583_),
    .A2(_03514_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08950_ (.A1(_03576_),
    .A2(_03571_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08951_ (.A1(_03563_),
    .A2(_03564_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08952_ (.A1(_03556_),
    .A2(_03552_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08953_ (.A1(_03536_),
    .A2(_03537_),
    .B(_03534_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _08954_ (.I(\as2650.debug_psl[3] ),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08955_ (.A1(_01516_),
    .A2(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08956_ (.A1(_03592_),
    .A2(_03594_),
    .B(_03538_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08957_ (.A1(_03550_),
    .A2(_03553_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08958_ (.A1(_03591_),
    .A2(_03595_),
    .B(_03596_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08959_ (.I(_03563_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08960_ (.A1(_03569_),
    .A2(_03571_),
    .B1(_03590_),
    .B2(_03597_),
    .C(_03598_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08961_ (.A1(_03528_),
    .A2(_03532_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08962_ (.A1(_03528_),
    .A2(_03531_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08963_ (.A1(_03600_),
    .A2(_03601_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _08964_ (.A1(_03589_),
    .A2(_03599_),
    .A3(_03602_),
    .B(_03600_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08965_ (.I(_03524_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08966_ (.A1(_03525_),
    .A2(_03603_),
    .B(_03604_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08967_ (.A1(_03583_),
    .A2(_03514_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08968_ (.A1(_03588_),
    .A2(_03605_),
    .B(_03606_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08969_ (.I(_03607_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08970_ (.A1(_01425_),
    .A2(_03505_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08971_ (.A1(_03506_),
    .A2(_03608_),
    .B(_03609_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08972_ (.A1(_03499_),
    .A2(_03587_),
    .A3(_03610_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08973_ (.A1(_01517_),
    .A2(_03499_),
    .B(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08974_ (.I(\as2650.debug_psl[0] ),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08975_ (.I(_03613_),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08976_ (.I(_01534_),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08977_ (.A1(_02152_),
    .A2(_02155_),
    .A3(_02157_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08978_ (.I(_03616_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08979_ (.I(_02257_),
    .Z(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08980_ (.A1(_03618_),
    .A2(_02930_),
    .A3(_02644_),
    .A4(_02161_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08981_ (.A1(_01160_),
    .A2(_01162_),
    .A3(_01317_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08982_ (.I(_01300_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08983_ (.A1(_01566_),
    .A2(_03619_),
    .B1(_03620_),
    .B2(_03621_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08984_ (.A1(_01792_),
    .A2(_03622_),
    .B(_03617_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08985_ (.I(_03519_),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08986_ (.A1(_03624_),
    .A2(_03498_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08987_ (.I(_03625_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08988_ (.A1(_03612_),
    .A2(_03626_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08989_ (.A1(_01225_),
    .A2(_03624_),
    .A3(_02285_),
    .A4(_01238_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08990_ (.I(_03628_),
    .Z(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08991_ (.I(_03629_),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08992_ (.A1(_01215_),
    .A2(_01301_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08993_ (.I(_03631_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08994_ (.I(_03632_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08995_ (.A1(_03630_),
    .A2(_03633_),
    .B(_01791_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08996_ (.A1(_03618_),
    .A2(_02162_),
    .A3(_02165_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08997_ (.I(_03635_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08998_ (.A1(_01148_),
    .A2(_01433_),
    .A3(_03496_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08999_ (.A1(_02156_),
    .A2(_03637_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09000_ (.A1(_03636_),
    .A2(_03004_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09001_ (.A1(_03614_),
    .A2(_03636_),
    .B(_03638_),
    .C(_03639_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09002_ (.A1(_03627_),
    .A2(_03634_),
    .A3(_03640_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09003_ (.A1(_01468_),
    .A2(_03617_),
    .B1(_03623_),
    .B2(_03641_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09004_ (.A1(_02667_),
    .A2(_03642_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09005_ (.A1(_03614_),
    .A2(_03615_),
    .B(_03643_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09006_ (.A1(_03493_),
    .A2(_03498_),
    .B1(_03644_),
    .B2(_01437_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09007_ (.I(_02163_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09008_ (.I(_02288_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09009_ (.A1(_03646_),
    .A2(_03647_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09010_ (.I(_02269_),
    .Z(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09011_ (.A1(_03649_),
    .A2(_03644_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09012_ (.I(_01424_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09013_ (.I(_03647_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09014_ (.A1(_03614_),
    .A2(_02352_),
    .B(_03649_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09015_ (.A1(_03651_),
    .A2(_03652_),
    .A3(_03653_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09016_ (.I(_03637_),
    .Z(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09017_ (.I(_03655_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09018_ (.A1(_03651_),
    .A2(_02289_),
    .B1(_03656_),
    .B2(_03612_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09019_ (.A1(_03656_),
    .A2(_03644_),
    .B(_03657_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09020_ (.A1(_03650_),
    .A2(_03654_),
    .B(_03658_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09021_ (.A1(_01518_),
    .A2(_02933_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09022_ (.A1(_02347_),
    .A2(_03660_),
    .B(_03650_),
    .C(_03648_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09023_ (.A1(_01237_),
    .A2(_01234_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09024_ (.I(_03662_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09025_ (.I(_03663_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09026_ (.A1(_03646_),
    .A2(_02271_),
    .A3(_03664_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09027_ (.A1(_01653_),
    .A2(_01435_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09028_ (.A1(_03665_),
    .A2(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09029_ (.A1(_03648_),
    .A2(_03659_),
    .B(_03661_),
    .C(_03667_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09030_ (.A1(_03493_),
    .A2(_03498_),
    .A3(_03612_),
    .B1(_03645_),
    .B2(_03668_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09031_ (.A1(_03491_),
    .A2(_03669_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09032_ (.A1(_03649_),
    .A2(_03665_),
    .A3(_01435_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(_02309_),
    .A2(_03651_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09034_ (.A1(_01760_),
    .A2(_02310_),
    .B(_03652_),
    .C(_03671_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09035_ (.A1(_02269_),
    .A2(_03647_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09036_ (.A1(_01191_),
    .A2(_01650_),
    .A3(_03673_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09037_ (.I(_03636_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09038_ (.I(_03617_),
    .Z(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09039_ (.A1(_03675_),
    .A2(_03676_),
    .B(_02173_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09040_ (.I(_02168_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09041_ (.A1(_02164_),
    .A2(_02158_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09042_ (.I(_03679_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09043_ (.A1(_03678_),
    .A2(_03063_),
    .B1(_03680_),
    .B2(net199),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09044_ (.A1(_01760_),
    .A2(_03677_),
    .B1(_03681_),
    .B2(_01152_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09045_ (.A1(_01651_),
    .A2(_03670_),
    .A3(_03672_),
    .B1(_03674_),
    .B2(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09046_ (.A1(_03491_),
    .A2(_03683_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09047_ (.A1(_03499_),
    .A2(_03656_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09048_ (.A1(_03507_),
    .A2(_03585_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09049_ (.A1(_03507_),
    .A2(_03607_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09050_ (.A1(_01236_),
    .A2(_01256_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09051_ (.I(_03687_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09052_ (.A1(_02643_),
    .A2(_01426_),
    .A3(_03687_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09053_ (.I(_03689_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09054_ (.A1(_02286_),
    .A2(_03506_),
    .A3(_03609_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09055_ (.A1(_03507_),
    .A2(_03688_),
    .B(_03690_),
    .C(_03691_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09056_ (.A1(_02155_),
    .A2(_03686_),
    .B(_03692_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09057_ (.A1(_03664_),
    .A2(_03685_),
    .B(_03693_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09058_ (.A1(_01209_),
    .A2(_01368_),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09059_ (.A1(_02285_),
    .A2(_01234_),
    .A3(_03695_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09060_ (.I(_03696_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09061_ (.A1(_03502_),
    .A2(_03697_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09062_ (.A1(_03694_),
    .A2(_03698_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _09063_ (.I(_03699_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09064_ (.A1(_01235_),
    .A2(_03498_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09065_ (.A1(_03506_),
    .A2(_03694_),
    .B1(_03700_),
    .B2(_03505_),
    .C(_03701_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09066_ (.I(_03495_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09067_ (.A1(_02930_),
    .A2(_03703_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09068_ (.A1(_03499_),
    .A2(_03626_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09069_ (.A1(_02168_),
    .A2(_03105_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09070_ (.A1(\as2650.debug_psl[2] ),
    .A2(_03636_),
    .B(_03705_),
    .C(_03706_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09071_ (.A1(_03702_),
    .A2(_03704_),
    .B(_03707_),
    .C(_03679_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09072_ (.A1(net210),
    .A2(_03680_),
    .B(_03708_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09073_ (.A1(_02667_),
    .A2(_03709_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09074_ (.A1(_01769_),
    .A2(_03615_),
    .B(_03710_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09075_ (.A1(_03701_),
    .A2(_03711_),
    .B(_03702_),
    .C(_02273_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09076_ (.A1(_02284_),
    .A2(_03712_),
    .B(_03667_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09077_ (.I(_03647_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09078_ (.A1(_01769_),
    .A2(_02323_),
    .B(_02373_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09079_ (.A1(_03714_),
    .A2(_03715_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09080_ (.A1(_01770_),
    .A2(_02284_),
    .A3(_02323_),
    .A4(_03648_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09081_ (.A1(_03712_),
    .A2(_03716_),
    .B(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09082_ (.A1(_03711_),
    .A2(_03713_),
    .B1(_03718_),
    .B2(_03667_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09083_ (.A1(_03493_),
    .A2(_03684_),
    .B(_03719_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09084_ (.A1(_03493_),
    .A2(_03702_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09085_ (.I(_01201_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09086_ (.A1(_03720_),
    .A2(_03721_),
    .B(_03722_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09087_ (.A1(_03651_),
    .A2(_02329_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09088_ (.A1(_03593_),
    .A2(_02330_),
    .B(_03652_),
    .C(_03723_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09089_ (.A1(_03678_),
    .A2(_03142_),
    .B1(_03680_),
    .B2(net214),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09090_ (.A1(_03593_),
    .A2(_03677_),
    .B1(_03725_),
    .B2(_01152_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09091_ (.A1(_01651_),
    .A2(_03670_),
    .A3(_03724_),
    .B1(_03726_),
    .B2(_03674_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09092_ (.A1(_03491_),
    .A2(_03727_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09093_ (.I(_01436_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09094_ (.A1(_02291_),
    .A2(_02449_),
    .B(_03714_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09095_ (.I(_00691_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09096_ (.I(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09097_ (.I(_03731_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09098_ (.A1(_03732_),
    .A2(_02338_),
    .B(_03665_),
    .C(_03649_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09099_ (.A1(_03233_),
    .A2(_03186_),
    .B(_03675_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09100_ (.I(_01802_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09101_ (.A1(_03735_),
    .A2(_03678_),
    .B(_03676_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09102_ (.A1(net215),
    .A2(_03233_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09103_ (.A1(_03732_),
    .A2(_02299_),
    .B1(_03734_),
    .B2(_03736_),
    .C1(_03737_),
    .C2(_03676_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09104_ (.A1(_03728_),
    .A2(_03729_),
    .A3(_03733_),
    .B1(_03674_),
    .B2(_03738_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09105_ (.A1(_03491_),
    .A2(_03739_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09106_ (.A1(_03492_),
    .A2(_03684_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09107_ (.A1(_03532_),
    .A2(_03697_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09108_ (.A1(_03574_),
    .A2(_03577_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09109_ (.I(_03602_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09110_ (.A1(_03742_),
    .A2(_03743_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09111_ (.I(_02154_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09112_ (.A1(_03589_),
    .A2(_03599_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09113_ (.A1(_03746_),
    .A2(_03743_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09114_ (.A1(_02287_),
    .A2(_03600_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09115_ (.A1(_02644_),
    .A2(_03601_),
    .A3(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09116_ (.A1(_03743_),
    .A2(_03695_),
    .B(_03696_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09117_ (.I(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09118_ (.A1(_03745_),
    .A2(_03747_),
    .B(_03749_),
    .C(_03751_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09119_ (.A1(_03663_),
    .A2(_03744_),
    .B(_03752_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09120_ (.A1(_03741_),
    .A2(_03753_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09121_ (.A1(_03664_),
    .A2(_03743_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09122_ (.A1(_03754_),
    .A2(_03755_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09123_ (.A1(_01530_),
    .A2(_02282_),
    .B(_02292_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09124_ (.A1(_03684_),
    .A2(_03756_),
    .B1(_03757_),
    .B2(_03673_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09125_ (.A1(_03673_),
    .A2(_03684_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09126_ (.A1(_02168_),
    .A2(_03223_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09127_ (.A1(_01529_),
    .A2(_03675_),
    .B(_03705_),
    .C(_03760_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09128_ (.A1(_03705_),
    .A2(_03756_),
    .B(_03761_),
    .C(_03634_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09129_ (.I(_01312_),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09130_ (.A1(_03763_),
    .A2(_03619_),
    .B1(_03620_),
    .B2(_01330_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09131_ (.A1(_01792_),
    .A2(_03764_),
    .B(_03617_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09132_ (.A1(net216),
    .A2(_03676_),
    .B1(_03762_),
    .B2(_03765_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09133_ (.A1(_02942_),
    .A2(_03766_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09134_ (.A1(_01530_),
    .A2(_02942_),
    .B(_03767_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09135_ (.A1(_01437_),
    .A2(_03759_),
    .B(_03768_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09136_ (.A1(_01437_),
    .A2(_03758_),
    .B(_03769_),
    .C(_03740_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09137_ (.A1(_03740_),
    .A2(_03756_),
    .B(_03770_),
    .C(_03303_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09138_ (.A1(\as2650.cycle[10] ),
    .A2(_01115_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09139_ (.I0(net8),
    .I1(net16),
    .I2(net32),
    .I3(net24),
    .S0(_01494_),
    .S1(_01496_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09140_ (.A1(_03771_),
    .A2(_03772_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09141_ (.I(\as2650.ext_io_addr[7] ),
    .Z(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _09142_ (.I0(net6),
    .I1(net30),
    .I2(net14),
    .I3(net22),
    .S0(\as2650.ext_io_addr[6] ),
    .S1(_03774_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09143_ (.I0(net3),
    .I1(net11),
    .I2(net27),
    .I3(net19),
    .S0(_03774_),
    .S1(_01496_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09144_ (.I(\as2650.ext_io_addr[6] ),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09145_ (.I0(net5),
    .I1(net13),
    .I2(net29),
    .I3(net21),
    .S0(_03774_),
    .S1(_03777_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09146_ (.A1(_03775_),
    .A2(_03776_),
    .A3(_03778_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09147_ (.I0(net7),
    .I1(net31),
    .I2(net15),
    .I3(net23),
    .S0(_03777_),
    .S1(_01494_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09148_ (.I0(net2),
    .I1(net26),
    .I2(net10),
    .I3(net18),
    .S0(\as2650.ext_io_addr[6] ),
    .S1(_03774_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09149_ (.I0(net4),
    .I1(net28),
    .I2(net12),
    .I3(net20),
    .S0(_03777_),
    .S1(_01494_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09150_ (.I0(net1),
    .I1(net9),
    .I2(net25),
    .I3(net17),
    .S0(\as2650.ext_io_addr[7] ),
    .S1(_03777_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09151_ (.A1(_03780_),
    .A2(_03781_),
    .A3(_03782_),
    .A4(_03783_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09152_ (.A1(_03779_),
    .A2(_03784_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09153_ (.A1(_03773_),
    .A2(_03785_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09154_ (.A1(_03618_),
    .A2(_03494_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09155_ (.A1(_02508_),
    .A2(_01642_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09156_ (.A1(_01403_),
    .A2(_01642_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09157_ (.A1(_02486_),
    .A2(_01632_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09158_ (.A1(_02341_),
    .A2(_01620_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09159_ (.A1(_02302_),
    .A2(_01568_),
    .B1(_01579_),
    .B2(_02307_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09160_ (.A1(_02308_),
    .A2(_01579_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09161_ (.A1(_02321_),
    .A2(_01588_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09162_ (.A1(_03792_),
    .A2(_03793_),
    .B(_03794_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09163_ (.A1(_02322_),
    .A2(_01589_),
    .B1(_01597_),
    .B2(_02326_),
    .C(_03795_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09164_ (.A1(_02326_),
    .A2(_01598_),
    .B1(_01610_),
    .B2(_02337_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09165_ (.A1(_02336_),
    .A2(_01610_),
    .B1(_01620_),
    .B2(_02340_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09166_ (.A1(_03796_),
    .A2(_03797_),
    .B(_03798_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09167_ (.A1(_03791_),
    .A2(_03799_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09168_ (.A1(_02486_),
    .A2(_01632_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09169_ (.A1(_03790_),
    .A2(_03800_),
    .B(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09170_ (.A1(_01758_),
    .A2(_02508_),
    .A3(_01642_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09171_ (.A1(_01758_),
    .A2(_03788_),
    .B1(_03789_),
    .B2(_03802_),
    .C(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09172_ (.A1(_03787_),
    .A2(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09173_ (.A1(_02943_),
    .A2(_02157_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09174_ (.A1(\as2650.debug_psu[5] ),
    .A2(\as2650.debug_psu[4] ),
    .A3(net181),
    .A4(_02248_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09175_ (.A1(_01900_),
    .A2(_02268_),
    .A3(_03807_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09176_ (.A1(_01758_),
    .A2(\as2650.debug_psl[2] ),
    .A3(_01791_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09177_ (.A1(_00707_),
    .A2(_01520_),
    .A3(_03614_),
    .A4(_01528_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _09178_ (.I(_01525_),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09179_ (.A1(_03811_),
    .A2(_02164_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09180_ (.A1(_03809_),
    .A2(_03810_),
    .B(_03812_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09181_ (.A1(_02951_),
    .A2(_03680_),
    .B(_03806_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09182_ (.I(_00771_),
    .Z(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09183_ (.A1(_00876_),
    .A2(_03815_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09184_ (.I(_00795_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09185_ (.A1(_01015_),
    .A2(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09186_ (.A1(_00820_),
    .A2(_00818_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09187_ (.A1(_03818_),
    .A2(_03819_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09188_ (.A1(_03816_),
    .A2(_03820_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09189_ (.I(_01475_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09190_ (.A1(_00856_),
    .A2(_03822_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09191_ (.I(_00877_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09192_ (.I(_03824_),
    .Z(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09193_ (.I(_00697_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09194_ (.A1(_03825_),
    .A2(_01471_),
    .B1(_01462_),
    .B2(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09195_ (.A1(_03826_),
    .A2(_03824_),
    .A3(_01470_),
    .A4(_01462_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09196_ (.A1(_03823_),
    .A2(_03827_),
    .B(_03828_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09197_ (.A1(_00877_),
    .A2(_01475_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09198_ (.A1(_00697_),
    .A2(_01469_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09199_ (.A1(_00856_),
    .A2(_01481_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09200_ (.A1(_03830_),
    .A2(_03831_),
    .A3(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09201_ (.A1(_03829_),
    .A2(_03833_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09202_ (.A1(_03829_),
    .A2(_03833_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09203_ (.A1(_03821_),
    .A2(_03834_),
    .B(_03835_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09204_ (.A1(_00694_),
    .A2(_03815_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09205_ (.I(_03817_),
    .Z(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09206_ (.A1(_00875_),
    .A2(_03838_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09207_ (.A1(_01016_),
    .A2(_00998_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09208_ (.A1(_03837_),
    .A2(_03839_),
    .A3(_03840_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09209_ (.I(_03825_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09210_ (.I(_03822_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09211_ (.I(_01471_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09212_ (.A1(_03842_),
    .A2(_03843_),
    .B1(_03844_),
    .B2(_00698_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09213_ (.I(_00698_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09214_ (.A1(_03846_),
    .A2(_00878_),
    .A3(_03843_),
    .A4(_03844_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09215_ (.A1(_03832_),
    .A2(_03845_),
    .B(_03847_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09216_ (.A1(_00856_),
    .A2(_00817_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09217_ (.A1(_03824_),
    .A2(_01481_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09218_ (.A1(_03826_),
    .A2(_03822_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09219_ (.A1(_03849_),
    .A2(_03850_),
    .A3(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09220_ (.A1(_03848_),
    .A2(_03852_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09221_ (.A1(_03841_),
    .A2(_03853_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09222_ (.A1(_03836_),
    .A2(_03854_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09223_ (.A1(_01012_),
    .A2(net189),
    .A3(_03820_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09224_ (.A1(_03818_),
    .A2(_03819_),
    .B(_03856_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09225_ (.A1(_03836_),
    .A2(_03854_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09226_ (.A1(_03857_),
    .A2(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09227_ (.I(_03837_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09228_ (.A1(_03839_),
    .A2(_03840_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09229_ (.A1(_03839_),
    .A2(_03840_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09230_ (.A1(_03860_),
    .A2(_03861_),
    .B(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09231_ (.A1(_03848_),
    .A2(_03852_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09232_ (.A1(_03841_),
    .A2(_03853_),
    .B(_03864_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09233_ (.A1(_01011_),
    .A2(net191),
    .B1(net190),
    .B2(_00695_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09234_ (.A1(_00694_),
    .A2(_01011_),
    .A3(_00998_),
    .A4(_01000_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09235_ (.I(_03867_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09236_ (.A1(_03866_),
    .A2(_03868_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09237_ (.I(_01482_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09238_ (.A1(_03842_),
    .A2(_03870_),
    .B1(_01477_),
    .B2(_03846_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09239_ (.A1(_03846_),
    .A2(_03842_),
    .A3(_03870_),
    .A4(_03843_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09240_ (.A1(_03849_),
    .A2(_03871_),
    .B(_03872_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09241_ (.A1(_03825_),
    .A2(_00818_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09242_ (.A1(_03826_),
    .A2(_01482_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09243_ (.A1(_00857_),
    .A2(_01015_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09244_ (.A1(_03874_),
    .A2(_03875_),
    .A3(_03876_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09245_ (.A1(_03873_),
    .A2(_03877_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09246_ (.A1(_03869_),
    .A2(_03878_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09247_ (.A1(_03865_),
    .A2(_03879_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09248_ (.A1(_03863_),
    .A2(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09249_ (.A1(_03855_),
    .A2(_03859_),
    .B(_03881_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09250_ (.A1(_01008_),
    .A2(_01005_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09251_ (.A1(_00817_),
    .A2(_00771_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09252_ (.I(_00821_),
    .Z(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09253_ (.A1(_01000_),
    .A2(_01483_),
    .B1(_01477_),
    .B2(_03885_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09254_ (.A1(_03885_),
    .A2(_03838_),
    .A3(_03870_),
    .A4(_01477_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09255_ (.A1(_03884_),
    .A2(_03886_),
    .B(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09256_ (.A1(_01011_),
    .A2(_01002_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09257_ (.A1(_03888_),
    .A2(_03889_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09258_ (.A1(_03883_),
    .A2(_03890_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09259_ (.A1(_03825_),
    .A2(_00857_),
    .A3(_01471_),
    .A4(_01463_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(_03817_),
    .A2(_01481_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09261_ (.A1(_00821_),
    .A2(_03822_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09262_ (.A1(_03884_),
    .A2(_03893_),
    .A3(_03894_),
    .Z(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09263_ (.I(_01470_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09264_ (.A1(_00997_),
    .A2(_03896_),
    .B1(_01463_),
    .B2(_00878_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09265_ (.A1(_03892_),
    .A2(_03895_),
    .A3(_03897_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09266_ (.A1(_03842_),
    .A2(_00997_),
    .A3(_01472_),
    .A4(_01464_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09267_ (.A1(_03824_),
    .A2(_01470_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09268_ (.A1(_00697_),
    .A2(_01462_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09269_ (.A1(_03900_),
    .A2(_03901_),
    .A3(_03823_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09270_ (.A1(_01015_),
    .A2(_03815_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09271_ (.A1(_00818_),
    .A2(_03817_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09272_ (.I(_00820_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09273_ (.A1(_03905_),
    .A2(_03870_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09274_ (.A1(_03903_),
    .A2(_03904_),
    .A3(_03906_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09275_ (.A1(_03899_),
    .A2(_03902_),
    .A3(_03907_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09276_ (.A1(_03898_),
    .A2(_03908_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09277_ (.A1(_03898_),
    .A2(_03908_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09278_ (.A1(_03891_),
    .A2(_03909_),
    .B(_03910_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09279_ (.A1(_03899_),
    .A2(_03902_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09280_ (.A1(_03899_),
    .A2(_03902_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09281_ (.A1(_03907_),
    .A2(_03912_),
    .B(_03913_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09282_ (.A1(_03834_),
    .A2(_03821_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09283_ (.A1(_03904_),
    .A2(_03906_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09284_ (.A1(_03904_),
    .A2(_03906_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09285_ (.A1(_03903_),
    .A2(_03916_),
    .B(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09286_ (.A1(_00695_),
    .A2(_01003_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09287_ (.A1(_03918_),
    .A2(_03919_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09288_ (.A1(_03914_),
    .A2(_03915_),
    .A3(_03920_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09289_ (.A1(_03911_),
    .A2(_03921_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09290_ (.A1(_01013_),
    .A2(net220),
    .A3(_03888_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09291_ (.A1(_03883_),
    .A2(_03890_),
    .B(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09292_ (.A1(_03911_),
    .A2(_03921_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09293_ (.A1(_03924_),
    .A2(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09294_ (.A1(_03922_),
    .A2(_03926_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09295_ (.A1(_03918_),
    .A2(_03919_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09296_ (.I(_03920_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09297_ (.A1(_03914_),
    .A2(_03915_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09298_ (.A1(_03914_),
    .A2(_03915_),
    .Z(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09299_ (.A1(_03929_),
    .A2(_03930_),
    .B(_03931_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09300_ (.A1(_03857_),
    .A2(_03858_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09301_ (.A1(_03932_),
    .A2(_03933_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09302_ (.A1(_03928_),
    .A2(_03934_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09303_ (.A1(_03927_),
    .A2(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09304_ (.A1(_00997_),
    .A2(_01465_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09305_ (.A1(_01482_),
    .A2(_03815_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09306_ (.A1(_00999_),
    .A2(_01476_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09307_ (.A1(_03905_),
    .A2(_03896_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09308_ (.A1(_03938_),
    .A2(_03939_),
    .A3(_03940_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09309_ (.A1(_03937_),
    .A2(_03941_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09310_ (.A1(_01017_),
    .A2(_00729_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09311_ (.A1(_01001_),
    .A2(_03843_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09312_ (.A1(_03838_),
    .A2(_03844_),
    .B1(_01464_),
    .B2(_03885_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09313_ (.A1(_03885_),
    .A2(_03838_),
    .A3(_03844_),
    .A4(_01463_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09314_ (.A1(_03944_),
    .A2(_03945_),
    .B(_03946_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09315_ (.A1(_01019_),
    .A2(_01002_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09316_ (.A1(_03943_),
    .A2(_03947_),
    .A3(_03948_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09317_ (.A1(_03942_),
    .A2(_03949_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09318_ (.A1(_03937_),
    .A2(_03941_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09319_ (.A1(_03892_),
    .A2(_03897_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09320_ (.A1(_03952_),
    .A2(_03895_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09321_ (.A1(_00876_),
    .A2(_00729_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09322_ (.A1(_00999_),
    .A2(_01476_),
    .B1(_03896_),
    .B2(_03905_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09323_ (.A1(_03905_),
    .A2(_00999_),
    .A3(_01476_),
    .A4(_03896_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09324_ (.A1(_03938_),
    .A2(_03955_),
    .B(_03956_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09325_ (.A1(_01017_),
    .A2(_01002_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09326_ (.A1(_03954_),
    .A2(_03957_),
    .A3(_03958_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09327_ (.A1(_03951_),
    .A2(_03953_),
    .A3(_03959_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(_03950_),
    .A2(_03960_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09329_ (.I(_03961_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09330_ (.A1(_03947_),
    .A2(_03948_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09331_ (.A1(_03947_),
    .A2(_03948_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09332_ (.A1(_03943_),
    .A2(_03963_),
    .B(_03964_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09333_ (.A1(_03950_),
    .A2(_03960_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09334_ (.A1(_03965_),
    .A2(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09335_ (.I(_03959_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09336_ (.A1(_03951_),
    .A2(_03953_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09337_ (.A1(_03951_),
    .A2(_03953_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09338_ (.A1(_03968_),
    .A2(_03969_),
    .B(_03970_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09339_ (.A1(_03891_),
    .A2(_03909_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09340_ (.A1(_03957_),
    .A2(_03958_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09341_ (.A1(_03957_),
    .A2(_03958_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09342_ (.A1(_03954_),
    .A2(_03973_),
    .B(_03974_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09343_ (.A1(_03971_),
    .A2(_03972_),
    .A3(_03975_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09344_ (.A1(_03962_),
    .A2(_03967_),
    .B(_03976_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09345_ (.A1(_01019_),
    .A2(_01005_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09346_ (.A1(_01483_),
    .A2(_00748_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09347_ (.A1(_01000_),
    .A2(_01001_),
    .A3(_01472_),
    .A4(_01465_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09348_ (.A1(_03978_),
    .A2(_03979_),
    .A3(_03980_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09349_ (.A1(net190),
    .A2(_01472_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09350_ (.A1(_00998_),
    .A2(_01464_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09351_ (.A1(_03982_),
    .A2(_03983_),
    .A3(_03944_),
    .Z(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09352_ (.A1(_03981_),
    .A2(_03984_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09353_ (.A1(_01001_),
    .A2(_01473_),
    .B1(_01465_),
    .B2(net190),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09354_ (.A1(_03980_),
    .A2(_03986_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09355_ (.A1(_01478_),
    .A2(_01003_),
    .B1(_01006_),
    .B2(_01484_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09356_ (.I(_03988_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09357_ (.A1(_01483_),
    .A2(_01478_),
    .A3(_01003_),
    .A4(_01005_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09358_ (.A1(_03987_),
    .A2(_03989_),
    .B(_03990_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09359_ (.A1(_03985_),
    .A2(_03991_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09360_ (.I(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09361_ (.A1(_01478_),
    .A2(_01004_),
    .A3(_01473_),
    .A4(_01007_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09362_ (.A1(_01479_),
    .A2(_01004_),
    .A3(_01474_),
    .A4(_01007_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09363_ (.A1(net189),
    .A2(_01466_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09364_ (.A1(_01004_),
    .A2(_01473_),
    .B1(_01006_),
    .B2(_01479_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09365_ (.A1(_03995_),
    .A2(_03996_),
    .A3(_03997_),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09366_ (.A1(_03990_),
    .A2(_03988_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09367_ (.A1(_03987_),
    .A2(_03999_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09368_ (.A1(_03994_),
    .A2(_03998_),
    .B(_04000_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09369_ (.A1(net220),
    .A2(_01474_),
    .A3(net219),
    .A4(_01466_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09370_ (.A1(_03995_),
    .A2(_03997_),
    .B(_03996_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09371_ (.A1(_03998_),
    .A2(_04002_),
    .A3(_04003_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09372_ (.A1(_03996_),
    .A2(_03997_),
    .B(_03994_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09373_ (.A1(_03987_),
    .A2(_03999_),
    .A3(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09374_ (.A1(_04004_),
    .A2(_04006_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09375_ (.A1(_03985_),
    .A2(_03991_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09376_ (.A1(_04001_),
    .A2(_04007_),
    .B(_04008_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09377_ (.A1(_03979_),
    .A2(_03980_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09378_ (.A1(_01019_),
    .A2(_01007_),
    .A3(_04010_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09379_ (.A1(_03979_),
    .A2(_03980_),
    .B(_04011_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09380_ (.A1(_03981_),
    .A2(_03984_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09381_ (.A1(_03942_),
    .A2(_03949_),
    .A3(_04013_),
    .Z(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09382_ (.A1(_04014_),
    .A2(_04012_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09383_ (.A1(_03993_),
    .A2(_04009_),
    .B(_04015_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09384_ (.A1(_03942_),
    .A2(_03949_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09385_ (.A1(_03950_),
    .A2(_04013_),
    .A3(_04017_),
    .B1(_04012_),
    .B2(_04014_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09386_ (.A1(_03950_),
    .A2(_03960_),
    .A3(_03965_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09387_ (.A1(_04019_),
    .A2(_04018_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09388_ (.A1(_04018_),
    .A2(_04019_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09389_ (.A1(_04016_),
    .A2(_04020_),
    .B(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09390_ (.A1(_03962_),
    .A2(_03967_),
    .A3(_03976_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09391_ (.A1(_03977_),
    .A2(_04022_),
    .B(_04023_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09392_ (.A1(_03971_),
    .A2(_03972_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09393_ (.A1(_03971_),
    .A2(_03972_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09394_ (.A1(_03975_),
    .A2(_04025_),
    .B(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09395_ (.A1(_03925_),
    .A2(_03924_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09396_ (.A1(_04027_),
    .A2(_04028_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09397_ (.A1(_04027_),
    .A2(_04028_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09398_ (.A1(_03927_),
    .A2(_03935_),
    .B1(_04024_),
    .B2(_04029_),
    .C(_04030_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09399_ (.A1(_03855_),
    .A2(_03859_),
    .A3(_03881_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09400_ (.A1(_03882_),
    .A2(_04032_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09401_ (.A1(_03932_),
    .A2(_03933_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09402_ (.A1(_03928_),
    .A2(_03934_),
    .B(_04034_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09403_ (.A1(_04033_),
    .A2(_04035_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09404_ (.A1(_04033_),
    .A2(_04035_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09405_ (.A1(_03936_),
    .A2(_04031_),
    .A3(_04036_),
    .B(_04037_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09406_ (.A1(_03863_),
    .A2(_03880_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09407_ (.A1(_03865_),
    .A2(_03879_),
    .B(_04039_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09408_ (.I(_03877_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09409_ (.A1(_03873_),
    .A2(_04041_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09410_ (.A1(_03869_),
    .A2(_03878_),
    .B(_04042_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09411_ (.A1(_01008_),
    .A2(net191),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09412_ (.A1(_03874_),
    .A2(_03875_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09413_ (.A1(_03874_),
    .A2(_03875_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09414_ (.A1(_03876_),
    .A2(_04045_),
    .B(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09415_ (.A1(_03846_),
    .A2(net193),
    .A3(_01016_),
    .A4(_00819_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09416_ (.A1(net193),
    .A2(_01016_),
    .B1(_00819_),
    .B2(_00996_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09417_ (.A1(_04048_),
    .A2(_04049_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09418_ (.A1(_01012_),
    .A2(net192),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09419_ (.A1(_04050_),
    .A2(_04051_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09420_ (.A1(_04047_),
    .A2(_04052_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09421_ (.A1(_04044_),
    .A2(_04053_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09422_ (.A1(_04043_),
    .A2(_04054_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09423_ (.A1(_03867_),
    .A2(_04055_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09424_ (.A1(_04040_),
    .A2(_04056_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09425_ (.A1(_04050_),
    .A2(_04051_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09426_ (.A1(_04048_),
    .A2(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09427_ (.A1(_00996_),
    .A2(_01017_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09428_ (.A1(_02969_),
    .A2(_00874_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09429_ (.A1(_04060_),
    .A2(_04061_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09430_ (.A1(_01008_),
    .A2(net192),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09431_ (.A1(_04062_),
    .A2(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09432_ (.A1(_04059_),
    .A2(_04064_),
    .Z(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09433_ (.A1(_04047_),
    .A2(_04052_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09434_ (.A1(_01009_),
    .A2(net191),
    .A3(_04053_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09435_ (.A1(_04066_),
    .A2(_04067_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09436_ (.A1(_04065_),
    .A2(_04068_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09437_ (.A1(_04043_),
    .A2(_04054_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09438_ (.A1(_03868_),
    .A2(_04055_),
    .B(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09439_ (.A1(_04069_),
    .A2(_04071_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09440_ (.A1(_04057_),
    .A2(_04072_),
    .Z(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09441_ (.A1(_04040_),
    .A2(_04056_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09442_ (.A1(_04057_),
    .A2(_04074_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09443_ (.I(_04075_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09444_ (.A1(_03882_),
    .A2(_04038_),
    .B(_04073_),
    .C(_04076_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09445_ (.I(_04071_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09446_ (.A1(_04057_),
    .A2(_04072_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09447_ (.A1(_04069_),
    .A2(_04078_),
    .B(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09448_ (.A1(_04065_),
    .A2(_04068_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09449_ (.A1(net194),
    .A2(_01018_),
    .A3(_04061_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09450_ (.A1(_04062_),
    .A2(_04063_),
    .B(_04082_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09451_ (.A1(_00996_),
    .A2(_01012_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09452_ (.A1(_01009_),
    .A2(net193),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09453_ (.A1(_04084_),
    .A2(_04085_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09454_ (.A1(_04083_),
    .A2(_04086_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09455_ (.A1(_04081_),
    .A2(_04087_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09456_ (.I(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09457_ (.A1(_00699_),
    .A2(_00693_),
    .A3(_04061_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09458_ (.A1(_04083_),
    .A2(_04086_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09459_ (.A1(_04059_),
    .A2(_04064_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(_04092_),
    .A2(_04087_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09461_ (.A1(_04091_),
    .A2(_04093_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09462_ (.A1(_04090_),
    .A2(_04094_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09463_ (.A1(_04089_),
    .A2(_04095_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09464_ (.I(_04096_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09465_ (.A1(_04092_),
    .A2(_04081_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09466_ (.A1(_04087_),
    .A2(_04098_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09467_ (.A1(_04077_),
    .A2(_04080_),
    .B(_04097_),
    .C(_04099_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09468_ (.A1(_04089_),
    .A2(_04095_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09469_ (.A1(_04061_),
    .A2(_04094_),
    .B(net194),
    .C(_01010_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09470_ (.A1(_04101_),
    .A2(_04102_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09471_ (.A1(_04100_),
    .A2(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09472_ (.A1(_04077_),
    .A2(_04080_),
    .B(_04099_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09473_ (.A1(_04105_),
    .A2(_04096_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09474_ (.A1(_04099_),
    .A2(_04077_),
    .A3(_04080_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09475_ (.A1(_04105_),
    .A2(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09476_ (.A1(_03882_),
    .A2(net351),
    .B(_04076_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09477_ (.A1(_04109_),
    .A2(_04073_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09478_ (.A1(_04075_),
    .A2(_03882_),
    .A3(net352),
    .Z(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09479_ (.A1(_03936_),
    .A2(_04031_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09480_ (.A1(_04112_),
    .A2(_04036_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09481_ (.A1(_04024_),
    .A2(_04029_),
    .B(_04030_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09482_ (.A1(_03927_),
    .A2(_03935_),
    .A3(_04114_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09483_ (.A1(_04024_),
    .A2(_04029_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09484_ (.A1(_03962_),
    .A2(_03967_),
    .A3(_03976_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09485_ (.A1(_04117_),
    .A2(_03977_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09486_ (.A1(_04022_),
    .A2(_04118_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09487_ (.A1(_04016_),
    .A2(_04020_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09488_ (.A1(_03993_),
    .A2(_04009_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09489_ (.A1(_04121_),
    .A2(_04015_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09490_ (.A1(_04001_),
    .A2(_04007_),
    .Z(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09491_ (.A1(_04123_),
    .A2(_04008_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09492_ (.A1(_04004_),
    .A2(_04006_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09493_ (.A1(_03998_),
    .A2(_04003_),
    .B(_04002_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09494_ (.A1(_04004_),
    .A2(_04126_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09495_ (.A1(_01578_),
    .A2(_02956_),
    .B1(_03539_),
    .B2(_00749_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09496_ (.A1(net219),
    .A2(_01467_),
    .B(_04127_),
    .C(_04128_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09497_ (.A1(_04122_),
    .A2(_04124_),
    .A3(_04125_),
    .A4(_04129_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09498_ (.A1(_04116_),
    .A2(_04119_),
    .A3(_04120_),
    .A4(_04130_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09499_ (.A1(_04115_),
    .A2(_04131_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09500_ (.A1(_04111_),
    .A2(_04113_),
    .A3(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09501_ (.A1(_04106_),
    .A2(_04108_),
    .A3(_04110_),
    .A4(_04133_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09502_ (.A1(_01224_),
    .A2(_01104_),
    .A3(_02932_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09503_ (.I(_04135_),
    .Z(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09504_ (.A1(_04104_),
    .A2(_04134_),
    .B(_04136_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09505_ (.A1(\as2650.debug_psl[6] ),
    .A2(_02167_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09506_ (.A1(_01536_),
    .A2(_04135_),
    .Z(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09507_ (.A1(_03635_),
    .A2(_03257_),
    .B(_04139_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09508_ (.A1(_01214_),
    .A2(_01432_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09509_ (.I(_04141_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09510_ (.A1(_04138_),
    .A2(_04140_),
    .B(_04142_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09511_ (.A1(_04137_),
    .A2(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09512_ (.I(_01578_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09513_ (.A1(_01014_),
    .A2(net216),
    .A3(_01020_),
    .A4(_01468_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09514_ (.A1(_03575_),
    .A2(_01587_),
    .A3(_04145_),
    .A4(_04146_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09515_ (.A1(_02954_),
    .A2(_04142_),
    .A3(_04147_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09516_ (.A1(_04144_),
    .A2(_04148_),
    .B(_03626_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09517_ (.I(_03516_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09518_ (.A1(_04150_),
    .A2(_03605_),
    .B(_02155_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09519_ (.A1(_04150_),
    .A2(_03605_),
    .B(_04151_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09520_ (.A1(_04150_),
    .A2(_03582_),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09521_ (.A1(_02287_),
    .A2(_03606_),
    .B(_03588_),
    .C(_02286_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09522_ (.A1(_03690_),
    .A2(_04154_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09523_ (.A1(_04150_),
    .A2(_03695_),
    .B(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09524_ (.A1(_03664_),
    .A2(_04153_),
    .B(_04156_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09525_ (.A1(_03583_),
    .A2(_03697_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09526_ (.A1(_04152_),
    .A2(_04157_),
    .B(_04158_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09527_ (.A1(_03741_),
    .A2(_03753_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09528_ (.A1(_03526_),
    .A2(_03579_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09529_ (.A1(_03526_),
    .A2(_03603_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09530_ (.A1(_01421_),
    .A2(_03604_),
    .B(_03525_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09531_ (.A1(_03526_),
    .A2(_03688_),
    .B1(_03690_),
    .B2(_03521_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09532_ (.A1(_03745_),
    .A2(_04162_),
    .B1(_04163_),
    .B2(_02286_),
    .C(_04164_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09533_ (.A1(_03663_),
    .A2(_04161_),
    .B(_04165_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09534_ (.A1(_03573_),
    .A2(_03566_),
    .A3(_03567_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09535_ (.A1(_01428_),
    .A2(_03574_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09536_ (.A1(_03590_),
    .A2(_03597_),
    .B(_03598_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09537_ (.A1(_03573_),
    .A2(_04169_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09538_ (.A1(_03576_),
    .A2(_03571_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09539_ (.A1(_02153_),
    .A2(_04171_),
    .B(_03589_),
    .C(_01127_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09540_ (.A1(_03573_),
    .A2(_03687_),
    .B1(_03689_),
    .B2(_03576_),
    .C(_04172_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09541_ (.A1(_03745_),
    .A2(_04170_),
    .B(_04173_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09542_ (.A1(_04167_),
    .A2(_04168_),
    .B(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09543_ (.A1(_03565_),
    .A2(_03597_),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09544_ (.A1(_03745_),
    .A2(_04176_),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09545_ (.A1(_03565_),
    .A2(_03555_),
    .A3(_03558_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09546_ (.A1(_03662_),
    .A2(_03566_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09547_ (.A1(_01127_),
    .A2(_03563_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09548_ (.A1(_02272_),
    .A2(_03564_),
    .B1(_04180_),
    .B2(_02153_),
    .C(_03689_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09549_ (.A1(_03565_),
    .A2(_03695_),
    .B1(_04178_),
    .B2(_04179_),
    .C(_04181_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _09550_ (.A1(_03560_),
    .A2(_03697_),
    .B1(_04177_),
    .B2(_04182_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09551_ (.A1(_03554_),
    .A2(_03688_),
    .B1(_03690_),
    .B2(_03550_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09552_ (.A1(_01425_),
    .A2(_01235_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09553_ (.A1(_03591_),
    .A2(_03595_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09554_ (.A1(_03554_),
    .A2(_03546_),
    .A3(_03547_),
    .Z(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09555_ (.A1(_03555_),
    .A2(_04187_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09556_ (.A1(_03550_),
    .A2(_03553_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09557_ (.A1(_02287_),
    .A2(_03596_),
    .B(_04189_),
    .C(_02285_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09558_ (.A1(_04185_),
    .A2(_04186_),
    .B1(_04188_),
    .B2(_03663_),
    .C(_04190_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09559_ (.A1(_04184_),
    .A2(_04191_),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09560_ (.A1(_03538_),
    .A2(_03544_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09561_ (.A1(_04193_),
    .A2(_03594_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09562_ (.A1(_04193_),
    .A2(_03545_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09563_ (.A1(_01425_),
    .A2(_03538_),
    .B(_03592_),
    .C(_02644_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09564_ (.A1(_04193_),
    .A2(_03688_),
    .B1(_03689_),
    .B2(_03543_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09565_ (.A1(_01428_),
    .A2(_04195_),
    .B(_04196_),
    .C(_04197_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09566_ (.A1(_04185_),
    .A2(_04194_),
    .B(_04198_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09567_ (.A1(_04175_),
    .A2(_04183_),
    .A3(_04192_),
    .A4(_04199_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09568_ (.A1(_04160_),
    .A2(_04166_),
    .A3(_04200_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09569_ (.A1(_03694_),
    .A2(_03698_),
    .B1(_04159_),
    .B2(_04201_),
    .C(_03637_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09570_ (.A1(_03703_),
    .A2(_04202_),
    .B(_03624_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09571_ (.A1(_03624_),
    .A2(_03495_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(_01010_),
    .A2(_01637_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09573_ (.A1(_01639_),
    .A2(_01300_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09574_ (.A1(_01014_),
    .A2(_01625_),
    .B(_04205_),
    .C(_04206_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09575_ (.A1(_01018_),
    .A2(_01616_),
    .B1(_01020_),
    .B2(_01302_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09576_ (.A1(_01607_),
    .A2(_01330_),
    .B1(_03575_),
    .B2(_01303_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09577_ (.A1(_01578_),
    .A2(_01340_),
    .B1(_03539_),
    .B2(_01341_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09578_ (.A1(_04208_),
    .A2(_04209_),
    .A3(_04210_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09579_ (.A1(net217),
    .A2(_01625_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09580_ (.A1(_00855_),
    .A2(_01324_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09581_ (.A1(_01484_),
    .A2(_01346_),
    .B1(_01480_),
    .B2(_01351_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09582_ (.I(_01285_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09583_ (.A1(_04145_),
    .A2(_01340_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09584_ (.A1(_01587_),
    .A2(_04215_),
    .B1(_01467_),
    .B2(_01359_),
    .C(_04216_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09585_ (.A1(_04212_),
    .A2(_04213_),
    .A3(_04214_),
    .A4(_04217_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09586_ (.A1(_01480_),
    .A2(_01351_),
    .B1(_04216_),
    .B2(_04210_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09587_ (.A1(_04219_),
    .A2(_04214_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09588_ (.A1(_04209_),
    .A2(_04220_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09589_ (.A1(_04208_),
    .A2(_04221_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09590_ (.A1(_01014_),
    .A2(_01625_),
    .B1(_04213_),
    .B2(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09591_ (.A1(\as2650.debug_psl[1] ),
    .A2(_01010_),
    .A3(_01637_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09592_ (.A1(\as2650.debug_psl[1] ),
    .A2(_04206_),
    .B1(_04207_),
    .B2(_04223_),
    .C(_04224_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09593_ (.A1(_04207_),
    .A2(_04211_),
    .A3(_04218_),
    .B(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09594_ (.A1(_04204_),
    .A2(_04226_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09595_ (.A1(_04149_),
    .A2(_04203_),
    .B(_04227_),
    .C(_03619_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09596_ (.A1(_03613_),
    .A2(_01790_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09597_ (.A1(_01790_),
    .A2(_01558_),
    .B(_04229_),
    .C(_03629_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09598_ (.A1(_03620_),
    .A2(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09599_ (.A1(_01594_),
    .A2(_01585_),
    .A3(_01286_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09600_ (.A1(_03621_),
    .A2(_03632_),
    .A3(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09601_ (.A1(_01626_),
    .A2(_01618_),
    .A3(_01604_),
    .A4(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09602_ (.A1(_04231_),
    .A2(_04234_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09603_ (.I(_01637_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09604_ (.A1(_01790_),
    .A2(_04236_),
    .B(_01296_),
    .C(_04229_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09605_ (.A1(_01627_),
    .A2(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09606_ (.A1(_04228_),
    .A2(_04235_),
    .B1(_04238_),
    .B2(_03633_),
    .C(_03616_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09607_ (.A1(_03806_),
    .A2(_03808_),
    .A3(_03813_),
    .B1(_03814_),
    .B2(_04239_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09608_ (.A1(_01520_),
    .A2(_02667_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09609_ (.A1(_03615_),
    .A2(_04240_),
    .B(_04241_),
    .C(_03655_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09610_ (.A1(_01254_),
    .A2(_01347_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09611_ (.A1(_04202_),
    .A2(_04243_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09612_ (.I(_01324_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09613_ (.A1(_03763_),
    .A2(_02590_),
    .B1(_02281_),
    .B2(_04245_),
    .C1(_04215_),
    .C2(_02408_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09614_ (.I(_01340_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09615_ (.A1(_02380_),
    .A2(_04247_),
    .B1(_02728_),
    .B2(_03621_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09616_ (.A1(_02302_),
    .A2(_01559_),
    .B1(_02327_),
    .B2(_01595_),
    .C(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09617_ (.A1(_01330_),
    .A2(_02448_),
    .B(_04243_),
    .C(_04249_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09618_ (.A1(_04246_),
    .A2(_04250_),
    .B(_03787_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09619_ (.A1(_04242_),
    .A2(_04244_),
    .B(_04251_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09620_ (.A1(_03805_),
    .A2(_04252_),
    .B(_02289_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09621_ (.I(_02268_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09622_ (.A1(_03615_),
    .A2(_04240_),
    .B(_04241_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09623_ (.A1(_04254_),
    .A2(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09624_ (.A1(_03646_),
    .A2(_02718_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09625_ (.A1(_01521_),
    .A2(_02718_),
    .B(_04257_),
    .C(_02283_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09626_ (.A1(_02273_),
    .A2(_04256_),
    .A3(_04258_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09627_ (.A1(_04253_),
    .A2(_04259_),
    .B(_03665_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09628_ (.A1(\as2650.debug_psu[7] ),
    .A2(_02267_),
    .B(_03812_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09629_ (.I(_02217_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09630_ (.I(_02267_),
    .Z(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09631_ (.A1(_04262_),
    .A2(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09632_ (.A1(_01769_),
    .A2(_02269_),
    .B(_04264_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09633_ (.I(_01870_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09634_ (.I(_04266_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09635_ (.A1(_01792_),
    .A2(_02268_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09636_ (.A1(_04267_),
    .A2(_04263_),
    .B(_04268_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09637_ (.I0(net181),
    .I1(_01520_),
    .S(_02267_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09638_ (.A1(_02812_),
    .A2(_04269_),
    .B1(_04270_),
    .B2(_02590_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09639_ (.A1(_02508_),
    .A2(_04261_),
    .B1(_04265_),
    .B2(_02323_),
    .C(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09640_ (.A1(_01843_),
    .A2(_02283_),
    .B(_03660_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09641_ (.A1(_02352_),
    .A2(_04273_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09642_ (.A1(\as2650.debug_psu[5] ),
    .A2(_02283_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09643_ (.A1(_01529_),
    .A2(_04254_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09644_ (.A1(_02342_),
    .A2(_04275_),
    .A3(_04276_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09645_ (.A1(_01759_),
    .A2(_04263_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09646_ (.A1(_01853_),
    .A2(_04254_),
    .B(_04278_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09647_ (.A1(_00691_),
    .A2(_02933_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09648_ (.A1(\as2650.debug_psu[4] ),
    .A2(_02933_),
    .B(_04280_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09649_ (.A1(_02309_),
    .A2(_04279_),
    .B1(_04281_),
    .B2(_02337_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09650_ (.A1(_04272_),
    .A2(_04274_),
    .A3(_04277_),
    .A4(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09651_ (.A1(_01429_),
    .A2(_04283_),
    .B(_03728_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09652_ (.A1(_01434_),
    .A2(_03492_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09653_ (.A1(_03787_),
    .A2(_03656_),
    .B(_04285_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09654_ (.A1(_03666_),
    .A2(_04255_),
    .B(_04286_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09655_ (.A1(_04260_),
    .A2(_04284_),
    .B(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09656_ (.A1(_01231_),
    .A2(_01212_),
    .A3(_01215_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09657_ (.A1(_00977_),
    .A2(_04289_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09658_ (.A1(_03805_),
    .A2(_04202_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09659_ (.A1(_04285_),
    .A2(_04291_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09660_ (.A1(_04290_),
    .A2(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09661_ (.A1(_02488_),
    .A2(_02342_),
    .A3(_02338_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09662_ (.A1(_02309_),
    .A2(_02304_),
    .A3(_02329_),
    .A4(_02324_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09663_ (.A1(_04294_),
    .A2(_04295_),
    .B(_02509_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09664_ (.A1(_04288_),
    .A2(_04293_),
    .B1(_04296_),
    .B2(_04290_),
    .C(_03771_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09665_ (.A1(_03786_),
    .A2(_04297_),
    .B(_03722_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09666_ (.A1(\as2650.cycle[8] ),
    .A2(_04289_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09667_ (.A1(_01449_),
    .A2(_01501_),
    .B1(_04298_),
    .B2(_02509_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09668_ (.A1(_02322_),
    .A2(_01589_),
    .B1(_01598_),
    .B2(_02327_),
    .C(_03792_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09669_ (.A1(_03798_),
    .A2(_03789_),
    .A3(_04300_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09670_ (.A1(_02322_),
    .A2(_01589_),
    .B1(_01610_),
    .B2(_02337_),
    .C(_03793_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09671_ (.A1(_02485_),
    .A2(_01632_),
    .Z(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09672_ (.A1(_02328_),
    .A2(_01598_),
    .B(_03791_),
    .C(_04303_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09673_ (.A1(_02303_),
    .A2(_01568_),
    .B(_04302_),
    .C(_04304_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09674_ (.A1(_04301_),
    .A2(_04305_),
    .B(_03703_),
    .C(_03804_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09675_ (.I(_04306_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09676_ (.A1(_03655_),
    .A2(_03700_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09677_ (.A1(_04307_),
    .A2(_04308_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09678_ (.A1(_04285_),
    .A2(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09679_ (.A1(_02943_),
    .A2(_02157_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09680_ (.I(_04261_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09681_ (.A1(_04204_),
    .A2(_04225_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09682_ (.A1(_02167_),
    .A2(_03296_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09683_ (.A1(_03811_),
    .A2(_02167_),
    .B(_04139_),
    .C(_04314_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09684_ (.A1(_04136_),
    .A2(_04104_),
    .B(_04142_),
    .C(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09685_ (.A1(_01639_),
    .A2(_04142_),
    .B(_04316_),
    .C(_03625_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09686_ (.A1(_04204_),
    .A2(_04317_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09687_ (.A1(_03638_),
    .A2(_03694_),
    .A3(_03698_),
    .B(_04318_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09688_ (.A1(_04313_),
    .A2(_04319_),
    .B(_03630_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09689_ (.A1(_03763_),
    .A2(_03633_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09690_ (.A1(_04231_),
    .A2(_04320_),
    .B(_04321_),
    .C(_03679_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09691_ (.A1(_02954_),
    .A2(_03616_),
    .B(_04311_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09692_ (.A1(_04311_),
    .A2(_04312_),
    .B1(_04322_),
    .B2(_04323_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09693_ (.I0(_03811_),
    .I1(_04324_),
    .S(_01534_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09694_ (.A1(_03655_),
    .A2(_04325_),
    .B(_04308_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09695_ (.A1(_03703_),
    .A2(_04243_),
    .A3(_04326_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09696_ (.A1(_02289_),
    .A2(_04306_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09697_ (.A1(_03646_),
    .A2(_02728_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09698_ (.A1(_01525_),
    .A2(_02728_),
    .B(_03673_),
    .C(_04329_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09699_ (.A1(_04327_),
    .A2(_04328_),
    .B(_04330_),
    .C(_01429_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09700_ (.A1(_01423_),
    .A2(_03728_),
    .A3(_02274_),
    .B(_04325_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09701_ (.A1(_03728_),
    .A2(_04331_),
    .B(_04332_),
    .C(_04286_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09702_ (.A1(_04310_),
    .A2(_04333_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09703_ (.A1(_04290_),
    .A2(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09704_ (.A1(_04299_),
    .A2(_04335_),
    .B(_01081_),
    .C(_03773_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09705_ (.I(_02696_),
    .Z(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09706_ (.A1(_01231_),
    .A2(_01363_),
    .B(_01213_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09707_ (.I(_04337_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09708_ (.A1(_01844_),
    .A2(_04338_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09709_ (.A1(_02266_),
    .A2(_03227_),
    .A3(_04338_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09710_ (.A1(_02275_),
    .A2(_04340_),
    .Z(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09711_ (.A1(_01104_),
    .A2(_02943_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09712_ (.A1(_02166_),
    .A2(_02259_),
    .A3(_04342_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09713_ (.A1(_02232_),
    .A2(_04343_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09714_ (.A1(_02159_),
    .A2(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09715_ (.A1(net188),
    .A2(_02174_),
    .B(_04345_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09716_ (.A1(_02974_),
    .A2(_04346_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09717_ (.A1(_01844_),
    .A2(_02316_),
    .B(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09718_ (.A1(_01843_),
    .A2(_02346_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09719_ (.A1(_02291_),
    .A2(_02346_),
    .B(_02274_),
    .C(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09720_ (.A1(_03016_),
    .A2(_04339_),
    .B(_04350_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09721_ (.A1(_04341_),
    .A2(_04348_),
    .B1(_04351_),
    .B2(_01655_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09722_ (.A1(_02791_),
    .A2(_04338_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09723_ (.I(_04353_),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09724_ (.I(_04354_),
    .Z(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09725_ (.A1(_02840_),
    .A2(_04339_),
    .B1(_04352_),
    .B2(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09726_ (.A1(_04336_),
    .A2(_04356_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09727_ (.I(_03424_),
    .Z(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09728_ (.I(_01852_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09729_ (.I(_04358_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09730_ (.A1(_02166_),
    .A2(_02261_),
    .B(_04357_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09731_ (.I(_04342_),
    .Z(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09732_ (.I(_04361_),
    .Z(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09733_ (.A1(_02166_),
    .A2(_02259_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09734_ (.I(_04363_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09735_ (.A1(_04357_),
    .A2(_04362_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09736_ (.A1(_04359_),
    .A2(_04362_),
    .B(_04364_),
    .C(_04365_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09737_ (.A1(_02174_),
    .A2(_04360_),
    .A3(_04366_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09738_ (.A1(_04145_),
    .A2(_02160_),
    .B(_04367_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09739_ (.A1(_02668_),
    .A2(_04368_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09740_ (.A1(_04359_),
    .A2(_02669_),
    .B(_04341_),
    .C(_04369_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09741_ (.A1(_01407_),
    .A2(_04338_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09742_ (.A1(_04254_),
    .A2(_01191_),
    .A3(_01429_),
    .A4(_01434_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09743_ (.A1(_01853_),
    .A2(_02381_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09744_ (.A1(_03714_),
    .A2(_04372_),
    .A3(_03671_),
    .A4(_04373_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09745_ (.A1(_01400_),
    .A2(_04357_),
    .A3(_04371_),
    .B(_04374_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09746_ (.A1(_01655_),
    .A2(_04375_),
    .B(_04354_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09747_ (.A1(_04357_),
    .A2(_04355_),
    .B1(_04370_),
    .B2(_04376_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09748_ (.A1(_04336_),
    .A2(_04377_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09749_ (.A1(_01862_),
    .A2(_03133_),
    .Z(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09750_ (.I(_04378_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09751_ (.A1(_01399_),
    .A2(_04378_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09752_ (.I(_01862_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09753_ (.A1(_04361_),
    .A2(_04379_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09754_ (.A1(_04381_),
    .A2(_04362_),
    .B(_04363_),
    .C(_04382_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09755_ (.A1(_02878_),
    .A2(_04364_),
    .B(_04383_),
    .C(_02159_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09756_ (.A1(net210),
    .A2(_02160_),
    .B(_04384_),
    .C(_02668_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09757_ (.A1(_04262_),
    .A2(_02669_),
    .B1(_04341_),
    .B2(_04380_),
    .C(_04385_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09758_ (.A1(_01399_),
    .A2(_04371_),
    .A3(_04378_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09759_ (.A1(_02291_),
    .A2(_02409_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09760_ (.A1(_01863_),
    .A2(_02409_),
    .B(_02290_),
    .C(_04388_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09761_ (.A1(_04387_),
    .A2(_04389_),
    .B(_03018_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09762_ (.A1(_04386_),
    .A2(_04390_),
    .B(_04354_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09763_ (.A1(_04355_),
    .A2(_04379_),
    .B(_04391_),
    .C(_03303_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09764_ (.A1(_01862_),
    .A2(_03123_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09765_ (.A1(_04266_),
    .A2(_04392_),
    .Z(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09766_ (.I(_02174_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09767_ (.A1(_04361_),
    .A2(_04393_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09768_ (.A1(_04267_),
    .A2(_04362_),
    .B(_04364_),
    .C(_04395_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09769_ (.A1(_02892_),
    .A2(_04364_),
    .B(_04396_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09770_ (.A1(_02160_),
    .A2(_04397_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09771_ (.A1(net214),
    .A2(_04394_),
    .B(_04398_),
    .C(_02668_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09772_ (.A1(_04267_),
    .A2(_02669_),
    .B(_04341_),
    .C(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09773_ (.A1(_01871_),
    .A2(_02812_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09774_ (.A1(_03714_),
    .A2(_04372_),
    .A3(_03723_),
    .A4(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09775_ (.A1(_01400_),
    .A2(_04371_),
    .A3(_04393_),
    .B(_04402_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09776_ (.A1(_01655_),
    .A2(_04403_),
    .B(_04354_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09777_ (.A1(_04355_),
    .A2(_04393_),
    .B1(_04400_),
    .B2(_04404_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09778_ (.A1(_04336_),
    .A2(_04405_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09779_ (.A1(_03233_),
    .A2(_03477_),
    .B(_03675_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09780_ (.A1(_01879_),
    .A2(_03678_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09781_ (.A1(_04394_),
    .A2(_04406_),
    .A3(_04407_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09782_ (.A1(_02284_),
    .A2(_02158_),
    .A3(_03737_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09783_ (.A1(_01879_),
    .A2(_01152_),
    .B(_04408_),
    .C(_04409_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09784_ (.A1(_01879_),
    .A2(_02450_),
    .B(_03729_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09785_ (.A1(_02738_),
    .A2(_02522_),
    .A3(_04372_),
    .A4(_04411_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09786_ (.A1(_02276_),
    .A2(_04410_),
    .B(_04412_),
    .C(_03303_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09787_ (.A1(net217),
    .A2(_04394_),
    .B1(_02169_),
    .B2(_02893_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09788_ (.A1(_02318_),
    .A2(_04413_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09789_ (.A1(_01894_),
    .A2(_02172_),
    .B(_04414_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09790_ (.A1(_02739_),
    .A2(_03652_),
    .A3(_04372_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09791_ (.A1(_01894_),
    .A2(_02719_),
    .B(_04257_),
    .C(_04416_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09792_ (.A1(_02276_),
    .A2(_04415_),
    .B1(_04417_),
    .B2(_01448_),
    .C(_02332_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09793_ (.A1(net218),
    .A2(_04394_),
    .B1(_02169_),
    .B2(_02924_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09794_ (.A1(_02318_),
    .A2(_04418_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09795_ (.A1(net37),
    .A2(_02172_),
    .B(_04419_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09796_ (.A1(_01900_),
    .A2(_02729_),
    .B(_04329_),
    .C(_04416_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09797_ (.A1(_02276_),
    .A2(_04420_),
    .B1(_04421_),
    .B2(_01448_),
    .C(_02332_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09798_ (.I(_01485_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09799_ (.I0(\as2650.irqs_latch[1] ),
    .I1(net44),
    .S(_04422_),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09800_ (.I(_04423_),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09801_ (.I(_01485_),
    .Z(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09802_ (.A1(net45),
    .A2(_04424_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09803_ (.A1(_02401_),
    .A2(_00010_),
    .B(_04425_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09804_ (.A1(net46),
    .A2(_04424_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09805_ (.A1(_02424_),
    .A2(_00010_),
    .B(_04426_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09806_ (.I0(\as2650.irqs_latch[4] ),
    .I1(\as2650.trap ),
    .S(_04422_),
    .Z(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09807_ (.I(_04427_),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09808_ (.A1(net47),
    .A2(_04424_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09809_ (.A1(_02403_),
    .A2(_00010_),
    .B(_04428_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09810_ (.A1(net48),
    .A2(_04422_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09811_ (.A1(_02400_),
    .A2(_04424_),
    .B(_04429_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09812_ (.I0(\as2650.irqs_latch[7] ),
    .I1(net49),
    .S(_04422_),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09813_ (.I(_04430_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09814_ (.I(_02165_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09815_ (.A1(_02661_),
    .A2(_01240_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09816_ (.A1(_01104_),
    .A2(_02299_),
    .A3(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09817_ (.A1(_02335_),
    .A2(_04431_),
    .A3(_04432_),
    .B1(_04433_),
    .B2(\as2650.trap ),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09818_ (.A1(_04336_),
    .A2(_04434_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09819_ (.I(\as2650.cycle[1] ),
    .Z(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09820_ (.I(_04435_),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09821_ (.I(\as2650.cycle[1] ),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09822_ (.A1(_04437_),
    .A2(net147),
    .B(_02971_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09823_ (.A1(_04436_),
    .A2(_01559_),
    .B(_04438_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09824_ (.A1(_04437_),
    .A2(net148),
    .B(_02971_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09825_ (.A1(_04436_),
    .A2(_01576_),
    .B(_04439_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09826_ (.I(_02970_),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09827_ (.A1(_04437_),
    .A2(net149),
    .B(_04440_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09828_ (.A1(_04436_),
    .A2(_01586_),
    .B(_04441_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09829_ (.A1(_04437_),
    .A2(net150),
    .B(_04440_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09830_ (.A1(_04436_),
    .A2(_01595_),
    .B(_04442_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09831_ (.I(_04435_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09832_ (.I(\as2650.cycle[1] ),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09833_ (.A1(_04444_),
    .A2(net151),
    .B(_04440_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09834_ (.A1(_04443_),
    .A2(_01605_),
    .B(_04445_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09835_ (.A1(_04444_),
    .A2(net152),
    .B(_04440_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09836_ (.A1(_04443_),
    .A2(_01618_),
    .B(_04446_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09837_ (.I(_02970_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09838_ (.A1(_04444_),
    .A2(net153),
    .B(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09839_ (.A1(_04443_),
    .A2(_01627_),
    .B(_04448_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09840_ (.A1(_04444_),
    .A2(net154),
    .B(_04447_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09841_ (.A1(_04443_),
    .A2(_01638_),
    .B(_04449_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09842_ (.A1(_01248_),
    .A2(net146),
    .B(\as2650.cycle[7] ),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09843_ (.A1(_01449_),
    .A2(_02650_),
    .A3(_04450_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09844_ (.I(_01439_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09845_ (.A1(net140),
    .A2(_01440_),
    .B(_04447_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09846_ (.A1(_02347_),
    .A2(_04451_),
    .B(_04452_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09847_ (.A1(net141),
    .A2(_01440_),
    .B(_04447_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09848_ (.A1(_02381_),
    .A2(_04451_),
    .B(_04453_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09849_ (.I(_02970_),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09850_ (.A1(net142),
    .A2(_01440_),
    .B(_04454_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09851_ (.A1(_02409_),
    .A2(_04451_),
    .B(_04455_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09852_ (.I(_01438_),
    .Z(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09853_ (.A1(net143),
    .A2(_04456_),
    .B(_04454_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09854_ (.A1(_02812_),
    .A2(_04451_),
    .B(_04457_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09855_ (.I(_01439_),
    .Z(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09856_ (.A1(net144),
    .A2(_04456_),
    .B(_04454_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09857_ (.A1(_02450_),
    .A2(_04458_),
    .B(_04459_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09858_ (.A1(net145),
    .A2(_04456_),
    .B(_04454_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09859_ (.A1(_02282_),
    .A2(_04458_),
    .B(_04460_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09860_ (.A1(_01496_),
    .A2(_04456_),
    .B(_01443_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09861_ (.A1(_02719_),
    .A2(_04458_),
    .B(_04461_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09862_ (.A1(_01495_),
    .A2(_01439_),
    .B(_01443_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09863_ (.A1(_02729_),
    .A2(_04458_),
    .B(_04462_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09864_ (.A1(_04435_),
    .A2(_01501_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09865_ (.A1(\as2650.io_bus_we ),
    .A2(_04435_),
    .B(_04463_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09866_ (.A1(_01449_),
    .A2(_02650_),
    .A3(_04464_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09867_ (.I(_00986_),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09868_ (.A1(net235),
    .A2(_04465_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09869_ (.A1(_01570_),
    .A2(_04466_),
    .B(_03722_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09870_ (.A1(_00956_),
    .A2(net237),
    .B(_02149_),
    .C(_01581_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09871_ (.A1(net222),
    .A2(_04465_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09872_ (.A1(_01590_),
    .A2(_04467_),
    .B(_03722_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09873_ (.A1(net223),
    .A2(_04465_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09874_ (.A1(_02139_),
    .A2(_01599_),
    .A3(_04468_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09875_ (.A1(net224),
    .A2(_04465_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09876_ (.A1(_01611_),
    .A2(_04469_),
    .B(_02297_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09877_ (.A1(_00951_),
    .A2(net237),
    .B(_02149_),
    .C(_01621_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09878_ (.A1(net226),
    .A2(_00986_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09879_ (.A1(_01633_),
    .A2(_04470_),
    .B(_02297_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09880_ (.A1(_00971_),
    .A2(net237),
    .B(_02149_),
    .C(_01643_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09881_ (.A1(_00588_),
    .A2(_02312_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09882_ (.I(_04471_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09883_ (.A1(_02351_),
    .A2(_04472_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09884_ (.A1(_02373_),
    .A2(_01405_),
    .A3(_01416_),
    .A4(_01268_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09885_ (.A1(_01190_),
    .A2(_01407_),
    .A3(_02354_),
    .A4(_04337_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09886_ (.A1(_01408_),
    .A2(_04474_),
    .B(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09887_ (.A1(_01431_),
    .A2(_04476_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09888_ (.A1(_04353_),
    .A2(_04477_),
    .B(_01175_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09889_ (.I(_04478_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09890_ (.I(_04479_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09891_ (.I(_04480_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09892_ (.A1(_01177_),
    .A2(_00974_),
    .A3(_01062_),
    .A4(_01076_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09893_ (.I(_04482_),
    .Z(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09894_ (.I(_04483_),
    .Z(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09895_ (.A1(_02270_),
    .A2(_04342_),
    .A3(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09896_ (.I(_04485_),
    .Z(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09897_ (.I(_04486_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09898_ (.I(_04485_),
    .Z(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09899_ (.A1(net188),
    .A2(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09900_ (.I(_04479_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09901_ (.I(_04490_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09902_ (.A1(_01518_),
    .A2(_04487_),
    .B(_04489_),
    .C(_04491_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09903_ (.A1(_04473_),
    .A2(_04481_),
    .B(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09904_ (.I(_04493_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09905_ (.I(_01870_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09906_ (.A1(_04262_),
    .A2(_04495_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09907_ (.I(_04482_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09908_ (.I(_04497_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09909_ (.A1(_04342_),
    .A2(_04498_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09910_ (.A1(_04499_),
    .A2(_04478_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09911_ (.A1(_02851_),
    .A2(_04500_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09912_ (.A1(_01853_),
    .A2(_04501_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09913_ (.A1(_04496_),
    .A2(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09914_ (.I(_04503_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09915_ (.I(_04504_),
    .Z(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09916_ (.I(_04503_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09917_ (.I(_04506_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09918_ (.A1(\as2650.stack[5][0] ),
    .A2(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09919_ (.A1(_04494_),
    .A2(_04505_),
    .B(_04508_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09920_ (.I(_04480_),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09921_ (.I(_04471_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09922_ (.I(_04471_),
    .Z(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09923_ (.A1(_02386_),
    .A2(_04511_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09924_ (.A1(_03065_),
    .A2(_04510_),
    .B(_04512_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09925_ (.I(_04486_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09926_ (.A1(net199),
    .A2(_04514_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09927_ (.A1(_01760_),
    .A2(_04487_),
    .B(_04491_),
    .C(_04515_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09928_ (.A1(_04509_),
    .A2(_04513_),
    .B(_04516_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09929_ (.I(_04517_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09930_ (.A1(\as2650.stack[5][1] ),
    .A2(_04507_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09931_ (.A1(_04505_),
    .A2(_04518_),
    .B(_04519_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09932_ (.I(_04471_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09933_ (.I0(_02413_),
    .I1(_03079_),
    .S(_04520_),
    .Z(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09934_ (.I(_04490_),
    .Z(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09935_ (.A1(net210),
    .A2(_04514_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09936_ (.A1(_01770_),
    .A2(_04487_),
    .B(_04522_),
    .C(_04523_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09937_ (.A1(_04509_),
    .A2(_04521_),
    .B(_04524_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09938_ (.I(_04525_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09939_ (.A1(\as2650.stack[5][2] ),
    .A2(_04507_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09940_ (.A1(_04505_),
    .A2(_04526_),
    .B(_04527_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09941_ (.I(_04472_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09942_ (.A1(_02429_),
    .A2(_04510_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09943_ (.A1(_02433_),
    .A2(_04528_),
    .B(_04529_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09944_ (.A1(net214),
    .A2(_04514_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09945_ (.A1(_03593_),
    .A2(_04487_),
    .B(_04522_),
    .C(_04531_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09946_ (.A1(_04509_),
    .A2(_04530_),
    .B(_04532_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09947_ (.I(_04533_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09948_ (.A1(\as2650.stack[5][3] ),
    .A2(_04507_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09949_ (.A1(_04505_),
    .A2(_04534_),
    .B(_04535_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09950_ (.I(_04504_),
    .Z(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09951_ (.A1(_03162_),
    .A2(_04510_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09952_ (.A1(_02472_),
    .A2(_04528_),
    .B(_04537_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09953_ (.I(_03730_),
    .Z(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09954_ (.I(_04486_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09955_ (.A1(net215),
    .A2(_04514_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09956_ (.A1(_04539_),
    .A2(_04540_),
    .B(_04522_),
    .C(_04541_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09957_ (.A1(_04509_),
    .A2(_04538_),
    .B(_04542_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09958_ (.I(_04543_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09959_ (.I(_04506_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09960_ (.A1(\as2650.stack[5][4] ),
    .A2(_04545_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09961_ (.A1(_04536_),
    .A2(_04544_),
    .B(_04546_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09962_ (.I(_04480_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09963_ (.A1(_03200_),
    .A2(_04511_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09964_ (.A1(_02494_),
    .A2(_04528_),
    .B(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09965_ (.I(_04498_),
    .Z(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09966_ (.A1(_02660_),
    .A2(_04361_),
    .A3(_04550_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09967_ (.I(_04551_),
    .Z(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09968_ (.I(_04551_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09969_ (.A1(_01529_),
    .A2(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09970_ (.A1(_02949_),
    .A2(_04552_),
    .B(_04522_),
    .C(_04554_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09971_ (.A1(_04547_),
    .A2(_04549_),
    .B(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09972_ (.I(_04556_),
    .Z(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09973_ (.A1(\as2650.stack[5][5] ),
    .A2(_04545_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09974_ (.A1(_04536_),
    .A2(_04557_),
    .B(_04558_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09975_ (.I0(_03234_),
    .I1(_03232_),
    .S(_04520_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09976_ (.I(_04490_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09977_ (.A1(_01521_),
    .A2(_04553_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09978_ (.A1(_02951_),
    .A2(_04552_),
    .B(_04560_),
    .C(_04561_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09979_ (.A1(_04547_),
    .A2(_04559_),
    .B(_04562_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09980_ (.I(_04563_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09981_ (.A1(\as2650.stack[5][6] ),
    .A2(_04545_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09982_ (.A1(_04536_),
    .A2(_04564_),
    .B(_04565_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09983_ (.A1(_03271_),
    .A2(_04511_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09984_ (.A1(_02513_),
    .A2(_04528_),
    .B(_04566_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09985_ (.A1(net218),
    .A2(_04488_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09986_ (.A1(_03811_),
    .A2(_04540_),
    .B(_04560_),
    .C(_04568_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09987_ (.A1(_04547_),
    .A2(_04567_),
    .B(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09988_ (.I(_04570_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09989_ (.A1(\as2650.stack[5][7] ),
    .A2(_04545_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09990_ (.A1(_04536_),
    .A2(_04571_),
    .B(_04572_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09991_ (.I(_04504_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09992_ (.I0(_03304_),
    .I1(_03307_),
    .S(_04520_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09993_ (.I(_04551_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09994_ (.A1(_01844_),
    .A2(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09995_ (.A1(_02956_),
    .A2(_04552_),
    .B(_04560_),
    .C(_04576_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09996_ (.A1(_04547_),
    .A2(_04574_),
    .B(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09997_ (.I(_04578_),
    .Z(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09998_ (.I(_04506_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09999_ (.A1(\as2650.stack[5][8] ),
    .A2(_04580_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10000_ (.A1(_04573_),
    .A2(_04579_),
    .B(_04581_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10001_ (.I(_04480_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10002_ (.I0(_03347_),
    .I1(_03345_),
    .S(_04520_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10003_ (.A1(net220),
    .A2(_04488_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10004_ (.A1(_04359_),
    .A2(_04540_),
    .B(_04560_),
    .C(_04584_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10005_ (.A1(_04582_),
    .A2(_04583_),
    .B(_04585_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10006_ (.I(_04586_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10007_ (.A1(\as2650.stack[5][9] ),
    .A2(_04580_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10008_ (.A1(_04573_),
    .A2(_04587_),
    .B(_04588_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10009_ (.A1(_02558_),
    .A2(_04511_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10010_ (.A1(_02562_),
    .A2(_04510_),
    .B(_04589_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10011_ (.I(_04490_),
    .Z(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10012_ (.A1(net189),
    .A2(_04488_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10013_ (.A1(_04262_),
    .A2(_04540_),
    .B(_04591_),
    .C(_04592_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10014_ (.A1(_04582_),
    .A2(_04590_),
    .B(_04593_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10015_ (.I(_04594_),
    .Z(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10016_ (.A1(\as2650.stack[5][10] ),
    .A2(_04580_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10017_ (.A1(_04573_),
    .A2(_04595_),
    .B(_04596_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10018_ (.I0(_03417_),
    .I1(_03419_),
    .S(_04472_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10019_ (.A1(_01871_),
    .A2(_04575_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10020_ (.A1(_00796_),
    .A2(_04552_),
    .B(_04591_),
    .C(_04598_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10021_ (.A1(_04582_),
    .A2(_04597_),
    .B(_04599_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10022_ (.I(_04600_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10023_ (.A1(\as2650.stack[5][11] ),
    .A2(_04580_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10024_ (.A1(_04573_),
    .A2(_04601_),
    .B(_04602_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10025_ (.I(_04504_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10026_ (.I0(_02598_),
    .I1(_02596_),
    .S(_04472_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10027_ (.A1(\as2650.debug_psu[4] ),
    .A2(_04575_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10028_ (.A1(_00822_),
    .A2(_04553_),
    .B(_04591_),
    .C(_04605_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10029_ (.A1(_04582_),
    .A2(_04604_),
    .B(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10030_ (.I(_04607_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10031_ (.I(_04506_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10032_ (.A1(\as2650.stack[5][12] ),
    .A2(_04609_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10033_ (.A1(_04603_),
    .A2(_04608_),
    .B(_04610_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10034_ (.I(_04486_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10035_ (.A1(_01887_),
    .A2(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10036_ (.A1(_02967_),
    .A2(_04611_),
    .B(_04612_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10037_ (.A1(_02830_),
    .A2(_04491_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10038_ (.A1(_04481_),
    .A2(_04613_),
    .B(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10039_ (.I(_04615_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10040_ (.A1(\as2650.stack[5][13] ),
    .A2(_04609_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10041_ (.A1(_04603_),
    .A2(_04616_),
    .B(_04617_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10042_ (.A1(_01894_),
    .A2(_04611_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10043_ (.A1(_02969_),
    .A2(_04611_),
    .B(_04618_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10044_ (.A1(_00932_),
    .A2(_04491_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10045_ (.A1(_04481_),
    .A2(_04619_),
    .B(_04620_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10046_ (.I(_04621_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10047_ (.A1(\as2650.stack[5][14] ),
    .A2(_04609_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10048_ (.A1(_04603_),
    .A2(_04622_),
    .B(_04623_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10049_ (.A1(_01900_),
    .A2(_04575_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10050_ (.A1(_00699_),
    .A2(_04553_),
    .B(_04591_),
    .C(_04624_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10051_ (.A1(\as2650.page_reg[2] ),
    .A2(_04481_),
    .B(_04625_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10052_ (.I(_04626_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10053_ (.A1(\as2650.stack[5][15] ),
    .A2(_04609_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10054_ (.A1(_04603_),
    .A2(_04627_),
    .B(_04628_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10055_ (.A1(_04499_),
    .A2(_04479_),
    .B(_02886_),
    .C(_04358_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10056_ (.A1(_04496_),
    .A2(_04629_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10057_ (.I(_04630_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10058_ (.I(_04631_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10059_ (.I(_04630_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10060_ (.I(_04633_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10061_ (.A1(\as2650.stack[6][0] ),
    .A2(_04634_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10062_ (.A1(_04494_),
    .A2(_04632_),
    .B(_04635_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10063_ (.A1(\as2650.stack[6][1] ),
    .A2(_04634_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10064_ (.A1(_04518_),
    .A2(_04632_),
    .B(_04636_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10065_ (.A1(\as2650.stack[6][2] ),
    .A2(_04634_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10066_ (.A1(_04526_),
    .A2(_04632_),
    .B(_04637_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10067_ (.A1(\as2650.stack[6][3] ),
    .A2(_04634_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10068_ (.A1(_04534_),
    .A2(_04632_),
    .B(_04638_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10069_ (.I(_04631_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10070_ (.I(_04633_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10071_ (.A1(\as2650.stack[6][4] ),
    .A2(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10072_ (.A1(_04544_),
    .A2(_04639_),
    .B(_04641_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10073_ (.A1(\as2650.stack[6][5] ),
    .A2(_04640_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10074_ (.A1(_04557_),
    .A2(_04639_),
    .B(_04642_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10075_ (.A1(\as2650.stack[6][6] ),
    .A2(_04640_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10076_ (.A1(_04564_),
    .A2(_04639_),
    .B(_04643_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10077_ (.A1(\as2650.stack[6][7] ),
    .A2(_04640_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10078_ (.A1(_04571_),
    .A2(_04639_),
    .B(_04644_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10079_ (.I(_04631_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10080_ (.I(_04633_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10081_ (.A1(\as2650.stack[6][8] ),
    .A2(_04646_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10082_ (.A1(_04579_),
    .A2(_04645_),
    .B(_04647_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10083_ (.A1(\as2650.stack[6][9] ),
    .A2(_04646_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10084_ (.A1(_04587_),
    .A2(_04645_),
    .B(_04648_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10085_ (.A1(\as2650.stack[6][10] ),
    .A2(_04646_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10086_ (.A1(_04595_),
    .A2(_04645_),
    .B(_04649_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10087_ (.A1(\as2650.stack[6][11] ),
    .A2(_04646_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10088_ (.A1(_04601_),
    .A2(_04645_),
    .B(_04650_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10089_ (.I(_04631_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10090_ (.I(_04633_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10091_ (.A1(\as2650.stack[6][12] ),
    .A2(_04652_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10092_ (.A1(_04608_),
    .A2(_04651_),
    .B(_04653_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10093_ (.A1(\as2650.stack[6][13] ),
    .A2(_04652_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10094_ (.A1(_04616_),
    .A2(_04651_),
    .B(_04654_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10095_ (.A1(\as2650.stack[6][14] ),
    .A2(_04652_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10096_ (.A1(_04622_),
    .A2(_04651_),
    .B(_04655_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10097_ (.A1(\as2650.stack[6][15] ),
    .A2(_04652_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10098_ (.A1(_04627_),
    .A2(_04651_),
    .B(_04656_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10099_ (.A1(_04499_),
    .A2(_04479_),
    .B(_02249_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10100_ (.A1(_04496_),
    .A2(_04657_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10101_ (.I(_04658_),
    .Z(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10102_ (.I(_04659_),
    .Z(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10103_ (.I(_04658_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10104_ (.I(_04661_),
    .Z(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10105_ (.A1(\as2650.stack[4][0] ),
    .A2(_04662_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10106_ (.A1(_04494_),
    .A2(_04660_),
    .B(_04663_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10107_ (.A1(\as2650.stack[4][1] ),
    .A2(_04662_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10108_ (.A1(_04518_),
    .A2(_04660_),
    .B(_04664_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10109_ (.A1(\as2650.stack[4][2] ),
    .A2(_04662_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10110_ (.A1(_04526_),
    .A2(_04660_),
    .B(_04665_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10111_ (.A1(\as2650.stack[4][3] ),
    .A2(_04662_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10112_ (.A1(_04534_),
    .A2(_04660_),
    .B(_04666_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10113_ (.I(_04659_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10114_ (.I(_04661_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10115_ (.A1(\as2650.stack[4][4] ),
    .A2(_04668_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10116_ (.A1(_04544_),
    .A2(_04667_),
    .B(_04669_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10117_ (.A1(\as2650.stack[4][5] ),
    .A2(_04668_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10118_ (.A1(_04557_),
    .A2(_04667_),
    .B(_04670_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10119_ (.A1(\as2650.stack[4][6] ),
    .A2(_04668_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10120_ (.A1(_04564_),
    .A2(_04667_),
    .B(_04671_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10121_ (.A1(\as2650.stack[4][7] ),
    .A2(_04668_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10122_ (.A1(_04571_),
    .A2(_04667_),
    .B(_04672_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10123_ (.I(_04659_),
    .Z(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10124_ (.I(_04661_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10125_ (.A1(\as2650.stack[4][8] ),
    .A2(_04674_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10126_ (.A1(_04579_),
    .A2(_04673_),
    .B(_04675_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10127_ (.A1(\as2650.stack[4][9] ),
    .A2(_04674_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10128_ (.A1(_04587_),
    .A2(_04673_),
    .B(_04676_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10129_ (.A1(\as2650.stack[4][10] ),
    .A2(_04674_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10130_ (.A1(_04595_),
    .A2(_04673_),
    .B(_04677_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10131_ (.A1(\as2650.stack[4][11] ),
    .A2(_04674_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10132_ (.A1(_04601_),
    .A2(_04673_),
    .B(_04678_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10133_ (.I(_04659_),
    .Z(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10134_ (.I(_04661_),
    .Z(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10135_ (.A1(\as2650.stack[4][12] ),
    .A2(_04680_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10136_ (.A1(_04608_),
    .A2(_04679_),
    .B(_04681_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10137_ (.A1(\as2650.stack[4][13] ),
    .A2(_04680_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10138_ (.A1(_04616_),
    .A2(_04679_),
    .B(_04682_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(\as2650.stack[4][14] ),
    .A2(_04680_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10140_ (.A1(_04622_),
    .A2(_04679_),
    .B(_04683_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10141_ (.A1(\as2650.stack[4][15] ),
    .A2(_04680_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10142_ (.A1(_04627_),
    .A2(_04679_),
    .B(_04684_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10143_ (.A1(_04359_),
    .A2(_04501_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10144_ (.A1(_04496_),
    .A2(_04685_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10145_ (.I(_04686_),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10146_ (.I(_04687_),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10147_ (.I(_04686_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10148_ (.I(_04689_),
    .Z(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10149_ (.A1(\as2650.stack[7][0] ),
    .A2(_04690_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10150_ (.A1(_04494_),
    .A2(_04688_),
    .B(_04691_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10151_ (.A1(\as2650.stack[7][1] ),
    .A2(_04690_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10152_ (.A1(_04518_),
    .A2(_04688_),
    .B(_04692_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10153_ (.A1(\as2650.stack[7][2] ),
    .A2(_04690_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10154_ (.A1(_04526_),
    .A2(_04688_),
    .B(_04693_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10155_ (.A1(\as2650.stack[7][3] ),
    .A2(_04690_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10156_ (.A1(_04534_),
    .A2(_04688_),
    .B(_04694_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10157_ (.I(_04687_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10158_ (.I(_04689_),
    .Z(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10159_ (.A1(\as2650.stack[7][4] ),
    .A2(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10160_ (.A1(_04544_),
    .A2(_04695_),
    .B(_04697_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10161_ (.A1(\as2650.stack[7][5] ),
    .A2(_04696_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10162_ (.A1(_04557_),
    .A2(_04695_),
    .B(_04698_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10163_ (.A1(\as2650.stack[7][6] ),
    .A2(_04696_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10164_ (.A1(_04564_),
    .A2(_04695_),
    .B(_04699_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10165_ (.A1(\as2650.stack[7][7] ),
    .A2(_04696_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10166_ (.A1(_04571_),
    .A2(_04695_),
    .B(_04700_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10167_ (.I(_04687_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10168_ (.I(_04689_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10169_ (.A1(\as2650.stack[7][8] ),
    .A2(_04702_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10170_ (.A1(_04579_),
    .A2(_04701_),
    .B(_04703_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10171_ (.A1(\as2650.stack[7][9] ),
    .A2(_04702_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10172_ (.A1(_04587_),
    .A2(_04701_),
    .B(_04704_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10173_ (.A1(\as2650.stack[7][10] ),
    .A2(_04702_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10174_ (.A1(_04595_),
    .A2(_04701_),
    .B(_04705_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10175_ (.A1(\as2650.stack[7][11] ),
    .A2(_04702_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10176_ (.A1(_04601_),
    .A2(_04701_),
    .B(_04706_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10177_ (.I(_04687_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10178_ (.I(_04689_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10179_ (.A1(\as2650.stack[7][12] ),
    .A2(_04708_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10180_ (.A1(_04608_),
    .A2(_04707_),
    .B(_04709_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10181_ (.A1(\as2650.stack[7][13] ),
    .A2(_04708_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10182_ (.A1(_04616_),
    .A2(_04707_),
    .B(_04710_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10183_ (.A1(\as2650.stack[7][14] ),
    .A2(_04708_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10184_ (.A1(_04622_),
    .A2(_04707_),
    .B(_04711_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10185_ (.A1(\as2650.stack[7][15] ),
    .A2(_04708_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10186_ (.A1(_04627_),
    .A2(_04707_),
    .B(_04712_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10187_ (.I(_04493_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10188_ (.I(_02247_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10189_ (.A1(_04714_),
    .A2(_04685_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10190_ (.I(_04715_),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10191_ (.I(_04716_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10192_ (.I(_04715_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10193_ (.I(_04718_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10194_ (.A1(\as2650.stack[3][0] ),
    .A2(_04719_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10195_ (.A1(_04713_),
    .A2(_04717_),
    .B(_04720_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10196_ (.I(_04517_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10197_ (.A1(\as2650.stack[3][1] ),
    .A2(_04719_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10198_ (.A1(_04721_),
    .A2(_04717_),
    .B(_04722_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10199_ (.I(_04525_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10200_ (.A1(\as2650.stack[3][2] ),
    .A2(_04719_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10201_ (.A1(_04723_),
    .A2(_04717_),
    .B(_04724_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10202_ (.I(_04533_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10203_ (.A1(\as2650.stack[3][3] ),
    .A2(_04719_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10204_ (.A1(_04725_),
    .A2(_04717_),
    .B(_04726_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10205_ (.I(_04543_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10206_ (.I(_04716_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10207_ (.I(_04718_),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10208_ (.A1(\as2650.stack[3][4] ),
    .A2(_04729_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10209_ (.A1(_04727_),
    .A2(_04728_),
    .B(_04730_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10210_ (.I(_04556_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10211_ (.A1(\as2650.stack[3][5] ),
    .A2(_04729_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10212_ (.A1(_04731_),
    .A2(_04728_),
    .B(_04732_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10213_ (.I(_04563_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10214_ (.A1(\as2650.stack[3][6] ),
    .A2(_04729_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10215_ (.A1(_04733_),
    .A2(_04728_),
    .B(_04734_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10216_ (.I(_04570_),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10217_ (.A1(\as2650.stack[3][7] ),
    .A2(_04729_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10218_ (.A1(_04735_),
    .A2(_04728_),
    .B(_04736_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10219_ (.I(_04578_),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10220_ (.I(_04716_),
    .Z(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10221_ (.I(_04718_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10222_ (.A1(\as2650.stack[3][8] ),
    .A2(_04739_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10223_ (.A1(_04737_),
    .A2(_04738_),
    .B(_04740_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10224_ (.I(_04586_),
    .Z(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10225_ (.A1(\as2650.stack[3][9] ),
    .A2(_04739_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10226_ (.A1(_04741_),
    .A2(_04738_),
    .B(_04742_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10227_ (.I(_04594_),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10228_ (.A1(\as2650.stack[3][10] ),
    .A2(_04739_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10229_ (.A1(_04743_),
    .A2(_04738_),
    .B(_04744_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10230_ (.I(_04600_),
    .Z(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10231_ (.A1(\as2650.stack[3][11] ),
    .A2(_04739_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10232_ (.A1(_04745_),
    .A2(_04738_),
    .B(_04746_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10233_ (.I(_04607_),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10234_ (.I(_04716_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10235_ (.I(_04718_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10236_ (.A1(\as2650.stack[3][12] ),
    .A2(_04749_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10237_ (.A1(_04747_),
    .A2(_04748_),
    .B(_04750_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10238_ (.I(_04615_),
    .Z(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10239_ (.A1(\as2650.stack[3][13] ),
    .A2(_04749_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10240_ (.A1(_04751_),
    .A2(_04748_),
    .B(_04752_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10241_ (.I(_04621_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10242_ (.A1(\as2650.stack[3][14] ),
    .A2(_04749_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10243_ (.A1(_04753_),
    .A2(_04748_),
    .B(_04754_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10244_ (.I(_04626_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10245_ (.A1(\as2650.stack[3][15] ),
    .A2(_04749_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10246_ (.A1(_04755_),
    .A2(_04748_),
    .B(_04756_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10247_ (.A1(_01075_),
    .A2(_03492_),
    .A3(_03497_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10248_ (.I(_04757_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10249_ (.I(_04758_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10250_ (.I(_04759_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10251_ (.I(_03783_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10252_ (.A1(_01077_),
    .A2(_03771_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10253_ (.I(_04762_),
    .Z(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10254_ (.A1(_01233_),
    .A2(_01075_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10255_ (.A1(_02791_),
    .A2(_04764_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10256_ (.I(_04765_),
    .Z(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10257_ (.A1(_02932_),
    .A2(_02258_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10258_ (.I(_04767_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10259_ (.A1(_04768_),
    .A2(_04497_),
    .Z(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10260_ (.I(_04768_),
    .Z(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10261_ (.I(_04482_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10262_ (.A1(_01128_),
    .A2(_01075_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10263_ (.A1(_03519_),
    .A2(_03495_),
    .B(_04141_),
    .C(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10264_ (.A1(_00975_),
    .A2(_01063_),
    .A3(_04773_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10265_ (.A1(_04770_),
    .A2(_04771_),
    .B1(_04774_),
    .B2(_01468_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10266_ (.A1(_01224_),
    .A2(_01227_),
    .A3(_03494_),
    .A4(_04772_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _10267_ (.A1(_00973_),
    .A2(_01062_),
    .A3(_04776_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10268_ (.I(_04777_),
    .Z(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10269_ (.I(_04778_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10270_ (.A1(_00980_),
    .A2(_01173_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10271_ (.A1(_01262_),
    .A2(_04780_),
    .B(_04773_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10272_ (.I(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10273_ (.I(_04776_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10274_ (.A1(_01566_),
    .A2(_01315_),
    .Z(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10275_ (.A1(_00976_),
    .A2(_01064_),
    .A3(_04783_),
    .B(_04784_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10276_ (.A1(_01558_),
    .A2(_04779_),
    .B1(_04782_),
    .B2(_01170_),
    .C(_04785_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10277_ (.A1(_03629_),
    .A2(_04482_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10278_ (.I(_04787_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10279_ (.A1(_01559_),
    .A2(_04769_),
    .B1(_04775_),
    .B2(_04786_),
    .C(_04788_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10280_ (.A1(_03629_),
    .A2(_04771_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10281_ (.A1(_03631_),
    .A2(_04497_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10282_ (.I(_04791_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10283_ (.A1(_01576_),
    .A2(_04790_),
    .B(_04792_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10284_ (.A1(_03632_),
    .A2(_04483_),
    .Z(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10285_ (.A1(_01791_),
    .A2(_04236_),
    .B(_04229_),
    .C(_04794_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10286_ (.A1(_01175_),
    .A2(_01398_),
    .A3(_01430_),
    .A4(_03637_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10287_ (.I(_04796_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10288_ (.A1(_04789_),
    .A2(_04793_),
    .B(_04795_),
    .C(_04797_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10289_ (.I(_04764_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10290_ (.A1(_01649_),
    .A2(_02833_),
    .A3(_04799_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10291_ (.I(_04800_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10292_ (.I(_04796_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10293_ (.A1(_04199_),
    .A2(_04802_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10294_ (.A1(_04801_),
    .A2(_04803_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10295_ (.A1(_01431_),
    .A2(_03147_),
    .A3(_04764_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10296_ (.A1(_01175_),
    .A2(_02635_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10297_ (.I(_04806_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10298_ (.A1(_01360_),
    .A2(_04805_),
    .B(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10299_ (.A1(_04798_),
    .A2(_04804_),
    .B(_04808_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10300_ (.I(_04806_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10301_ (.A1(_02612_),
    .A2(_02633_),
    .B(_01251_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10302_ (.A1(_02646_),
    .A2(_04811_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10303_ (.I(_04812_),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10304_ (.A1(_01558_),
    .A2(_04813_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10305_ (.I(_04765_),
    .Z(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10306_ (.A1(_04810_),
    .A2(_04814_),
    .B(_04815_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10307_ (.A1(_01174_),
    .A2(_04298_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10308_ (.I(_04817_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10309_ (.A1(_01360_),
    .A2(_04766_),
    .B1(_04809_),
    .B2(_04816_),
    .C(_04818_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10310_ (.A1(_01076_),
    .A2(_04290_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10311_ (.I(_04820_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10312_ (.I(_04762_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10313_ (.A1(_02303_),
    .A2(_04821_),
    .B(_04822_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10314_ (.A1(_04761_),
    .A2(_04763_),
    .B1(_04819_),
    .B2(_04823_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10315_ (.I(_04758_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10316_ (.A1(_04199_),
    .A2(_04825_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10317_ (.A1(_04760_),
    .A2(_04824_),
    .B(_04826_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10318_ (.I(_04827_),
    .Z(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10319_ (.I(_04828_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10320_ (.A1(_04136_),
    .A2(_04498_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10321_ (.A1(_01251_),
    .A2(_02162_),
    .A3(_04431_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10322_ (.A1(_04831_),
    .A2(_04497_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10323_ (.I(_04832_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10324_ (.I(_04833_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10325_ (.A1(_01204_),
    .A2(_03618_),
    .A3(_01240_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10326_ (.A1(_01171_),
    .A2(_01077_),
    .A3(_04431_),
    .A4(_04835_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10327_ (.A1(_04830_),
    .A2(_04834_),
    .A3(_04836_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10328_ (.A1(_01629_),
    .A2(_04758_),
    .B(_02163_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10329_ (.I(_04838_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10330_ (.A1(_01629_),
    .A2(_04759_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10331_ (.A1(_02635_),
    .A2(_01174_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10332_ (.A1(_01178_),
    .A2(_04781_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10333_ (.A1(\as2650.cycle[10] ),
    .A2(_01115_),
    .A3(_01173_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10334_ (.A1(_04777_),
    .A2(_04842_),
    .A3(_04817_),
    .A4(_04843_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10335_ (.A1(_02370_),
    .A2(_04799_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10336_ (.A1(_04757_),
    .A2(_04841_),
    .A3(_04844_),
    .A4(_04845_),
    .Z(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10337_ (.A1(_01076_),
    .A2(_01190_),
    .A3(_01649_),
    .A4(_03497_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10338_ (.A1(_01363_),
    .A2(_01452_),
    .B(_01381_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10339_ (.A1(_04767_),
    .A2(_03628_),
    .A3(_03631_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10340_ (.A1(_01149_),
    .A2(_01174_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10341_ (.A1(_04848_),
    .A2(_04849_),
    .B(_04850_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _10342_ (.A1(_04846_),
    .A2(_04847_),
    .A3(_04851_),
    .A4(_04800_),
    .Z(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10343_ (.A1(_04263_),
    .A2(_04852_),
    .Z(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10344_ (.A1(_04840_),
    .A2(_04853_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10345_ (.A1(_03730_),
    .A2(_04839_),
    .A3(_04854_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10346_ (.A1(_04837_),
    .A2(_04855_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10347_ (.I(_04856_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10348_ (.I(_04830_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10349_ (.A1(_04116_),
    .A2(_04858_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10350_ (.A1(_04831_),
    .A2(_04484_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10351_ (.I(_04860_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10352_ (.I(_04861_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10353_ (.I(_04861_),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10354_ (.A1(_03539_),
    .A2(_04863_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10355_ (.A1(_04136_),
    .A2(_04484_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10356_ (.I(_04865_),
    .Z(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10357_ (.I(_04866_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10358_ (.A1(_03336_),
    .A2(_04862_),
    .B(_04864_),
    .C(_04867_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10359_ (.A1(_04859_),
    .A2(_04868_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10360_ (.A1(_03731_),
    .A2(_04837_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10361_ (.I(_04870_),
    .Z(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10362_ (.A1(_02572_),
    .A2(_04870_),
    .A3(_04855_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10363_ (.I(_04872_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10364_ (.A1(_04869_),
    .A2(_04871_),
    .B1(_04873_),
    .B2(\as2650.regs[5][0] ),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10365_ (.A1(_04829_),
    .A2(_04857_),
    .B(_04874_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10366_ (.I(_04759_),
    .Z(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10367_ (.I(_03781_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10368_ (.I(_04762_),
    .Z(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10369_ (.I(_04791_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10370_ (.I(_01358_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10371_ (.A1(_00975_),
    .A2(_01064_),
    .A3(_04783_),
    .B(_04879_),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10372_ (.A1(_01576_),
    .A2(_04779_),
    .B1(_04782_),
    .B2(_01169_),
    .C(_04880_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10373_ (.A1(_04768_),
    .A2(_04483_),
    .B1(_04774_),
    .B2(net199),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10374_ (.A1(_01528_),
    .A2(_04247_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10375_ (.A1(_04881_),
    .A2(_04882_),
    .B1(_04883_),
    .B2(_04769_),
    .C(_04787_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10376_ (.A1(_01586_),
    .A2(_04790_),
    .B(_04792_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10377_ (.A1(_01566_),
    .A2(_04878_),
    .B1(_04884_),
    .B2(_04885_),
    .C(_04797_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10378_ (.A1(_04192_),
    .A2(_04802_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10379_ (.A1(_04801_),
    .A2(_04887_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10380_ (.A1(_01358_),
    .A2(_04805_),
    .B(_04807_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10381_ (.A1(_04886_),
    .A2(_04888_),
    .B(_04889_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10382_ (.I(_04812_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10383_ (.A1(_02639_),
    .A2(_02623_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10384_ (.A1(_01356_),
    .A2(_04892_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(_04813_),
    .A2(_04893_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10386_ (.I(_04841_),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10387_ (.A1(_04247_),
    .A2(_04891_),
    .B(_04894_),
    .C(_04895_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10388_ (.A1(_04766_),
    .A2(_04896_),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10389_ (.I(_04818_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10390_ (.A1(_01358_),
    .A2(_04766_),
    .B1(_04890_),
    .B2(_04897_),
    .C(_04898_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10391_ (.A1(_02308_),
    .A2(_04821_),
    .B(_04763_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10392_ (.A1(_04876_),
    .A2(_04877_),
    .B1(_04899_),
    .B2(_04900_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10393_ (.A1(_04192_),
    .A2(_04825_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10394_ (.A1(_04875_),
    .A2(_04901_),
    .B(_04902_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10395_ (.I(_04903_),
    .Z(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10396_ (.I(_04904_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10397_ (.I(_04872_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10398_ (.I(_04830_),
    .Z(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10399_ (.I(_04907_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10400_ (.A1(_04115_),
    .A2(_04908_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10401_ (.I(_04861_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10402_ (.I(_04861_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10403_ (.A1(_04145_),
    .A2(_04911_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10404_ (.I(_04866_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10405_ (.A1(_03373_),
    .A2(_04910_),
    .B(_04912_),
    .C(_04913_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10406_ (.A1(_04909_),
    .A2(_04914_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10407_ (.I(_04870_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10408_ (.A1(\as2650.regs[5][1] ),
    .A2(_04906_),
    .B1(_04915_),
    .B2(_04916_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10409_ (.A1(_04857_),
    .A2(_04905_),
    .B(_04917_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10410_ (.I(_04183_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10411_ (.I(_04760_),
    .Z(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10412_ (.I(_04820_),
    .Z(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10413_ (.I(_04841_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10414_ (.I(_04847_),
    .Z(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10415_ (.A1(\as2650.debug_psl[5] ),
    .A2(_01286_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10416_ (.A1(_01585_),
    .A2(_04923_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10417_ (.A1(_04768_),
    .A2(_04483_),
    .B1(_04774_),
    .B2(_01480_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10418_ (.I(_01355_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10419_ (.A1(_00975_),
    .A2(_01063_),
    .A3(_04783_),
    .B(_04926_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10420_ (.A1(_01585_),
    .A2(_04778_),
    .B1(_04782_),
    .B2(_01169_),
    .C(_04927_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10421_ (.A1(_04769_),
    .A2(_04924_),
    .B1(_04925_),
    .B2(_04928_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10422_ (.A1(_01594_),
    .A2(_04788_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10423_ (.A1(_04788_),
    .A2(_04929_),
    .B(_04930_),
    .C(_04792_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10424_ (.A1(_04247_),
    .A2(_04794_),
    .B(_04922_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10425_ (.A1(_04183_),
    .A2(_04922_),
    .B1(_04931_),
    .B2(_04932_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10426_ (.I(_04812_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10427_ (.A1(_02613_),
    .A2(_02653_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10428_ (.A1(_01352_),
    .A2(_04935_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10429_ (.A1(_02639_),
    .A2(_01353_),
    .B(_04813_),
    .C(_04936_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10430_ (.A1(_01586_),
    .A2(_04934_),
    .B(_04937_),
    .C(_04895_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10431_ (.A1(_04921_),
    .A2(_04933_),
    .B(_04938_),
    .C(_04815_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10432_ (.I(_04845_),
    .Z(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10433_ (.A1(_01355_),
    .A2(_04940_),
    .B(_04920_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10434_ (.A1(_02408_),
    .A2(_04920_),
    .B1(_04939_),
    .B2(_04941_),
    .C(_04822_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10435_ (.A1(_03776_),
    .A2(_04877_),
    .B(_04942_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10436_ (.A1(_04875_),
    .A2(_04943_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10437_ (.A1(_04918_),
    .A2(_04919_),
    .B(_04944_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10438_ (.I(_04945_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10439_ (.A1(_01587_),
    .A2(_04863_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10440_ (.I(_04865_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10441_ (.I(_04948_),
    .Z(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10442_ (.A1(_03411_),
    .A2(_04862_),
    .B(_04947_),
    .C(_04949_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10443_ (.A1(_04113_),
    .A2(_04913_),
    .B(_04950_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10444_ (.A1(\as2650.regs[5][2] ),
    .A2(_04906_),
    .B1(_04951_),
    .B2(_04916_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10445_ (.A1(_04857_),
    .A2(_04946_),
    .B(_04952_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10446_ (.I(_03782_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10447_ (.I(_04778_),
    .Z(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10448_ (.A1(_00976_),
    .A2(_01064_),
    .A3(_04783_),
    .B(_01350_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10449_ (.A1(_01594_),
    .A2(_04954_),
    .B1(_04782_),
    .B2(_01170_),
    .C(_04955_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10450_ (.I(_04774_),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10451_ (.A1(_04770_),
    .A2(_04771_),
    .B1(_04957_),
    .B2(_01484_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10452_ (.A1(_04215_),
    .A2(_04923_),
    .B(_01528_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10453_ (.A1(_01346_),
    .A2(_04959_),
    .Z(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10454_ (.A1(_04956_),
    .A2(_04958_),
    .B1(_04960_),
    .B2(_04769_),
    .C(_04788_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10455_ (.A1(_01605_),
    .A2(_04790_),
    .B(_04878_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10456_ (.I(_04796_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10457_ (.A1(_04215_),
    .A2(_04878_),
    .B1(_04961_),
    .B2(_04962_),
    .C(_04963_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10458_ (.A1(_04175_),
    .A2(_04797_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10459_ (.A1(_04801_),
    .A2(_04965_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10460_ (.I(_01350_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10461_ (.A1(_04967_),
    .A2(_04805_),
    .B(_04810_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10462_ (.A1(_04964_),
    .A2(_04966_),
    .B(_04968_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10463_ (.I(_04892_),
    .Z(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10464_ (.A1(_02640_),
    .A2(_01348_),
    .B1(_04970_),
    .B2(_01344_),
    .C(_04934_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10465_ (.A1(_01303_),
    .A2(_04891_),
    .B(_04971_),
    .C(_04895_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10466_ (.A1(_04766_),
    .A2(_04972_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10467_ (.A1(_01350_),
    .A2(_04940_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10468_ (.A1(_04969_),
    .A2(_04973_),
    .B(_04974_),
    .C(_04898_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10469_ (.A1(_02328_),
    .A2(_04821_),
    .B(_04763_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10470_ (.A1(_04953_),
    .A2(_04877_),
    .B1(_04975_),
    .B2(_04976_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10471_ (.A1(_04175_),
    .A2(_04760_),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10472_ (.A1(_04875_),
    .A2(_04977_),
    .B(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10473_ (.I(_04979_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10474_ (.A1(_03575_),
    .A2(_04863_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10475_ (.A1(_03444_),
    .A2(_04862_),
    .B(_04981_),
    .C(_04949_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10476_ (.A1(_04111_),
    .A2(_04913_),
    .B(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10477_ (.A1(\as2650.regs[5][3] ),
    .A2(_04906_),
    .B1(_04983_),
    .B2(_04916_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10478_ (.A1(_04857_),
    .A2(_04980_),
    .B(_04984_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10479_ (.I(_04856_),
    .Z(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10480_ (.I(_01336_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10481_ (.I0(_01604_),
    .I1(_04986_),
    .S(_04778_),
    .Z(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10482_ (.A1(net215),
    .A2(_04957_),
    .B1(_04987_),
    .B2(_04842_),
    .C(_04787_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10483_ (.A1(_04245_),
    .A2(_04790_),
    .B(_04792_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10484_ (.A1(_01595_),
    .A2(_04878_),
    .B1(_04988_),
    .B2(_04989_),
    .C(_04802_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10485_ (.A1(_04160_),
    .A2(_04922_),
    .B(_04801_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10486_ (.A1(_01336_),
    .A2(_04805_),
    .B(_04807_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10487_ (.A1(_04990_),
    .A2(_04991_),
    .B(_04992_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10488_ (.A1(_02614_),
    .A2(_01334_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10489_ (.A1(_01331_),
    .A2(_04970_),
    .B(_04994_),
    .C(_04813_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10490_ (.A1(_01605_),
    .A2(_04934_),
    .B(_04995_),
    .C(_04895_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10491_ (.A1(_04815_),
    .A2(_04996_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10492_ (.A1(_04986_),
    .A2(_04845_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10493_ (.A1(_04993_),
    .A2(_04997_),
    .B(_04998_),
    .C(_04818_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10494_ (.A1(_02449_),
    .A2(_04920_),
    .B(_04822_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10495_ (.A1(_03778_),
    .A2(_04763_),
    .B1(_04999_),
    .B2(_05000_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10496_ (.I0(_05001_),
    .I1(_04160_),
    .S(_04759_),
    .Z(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10497_ (.I(_05002_),
    .Z(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10498_ (.I(_05003_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10499_ (.A1(_04110_),
    .A2(_04908_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10500_ (.A1(_01607_),
    .A2(_04911_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10501_ (.A1(_03477_),
    .A2(_04910_),
    .B(_05006_),
    .C(_04913_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10502_ (.A1(_05005_),
    .A2(_05007_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10503_ (.A1(\as2650.regs[5][4] ),
    .A2(_04906_),
    .B1(_05008_),
    .B2(_04916_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10504_ (.A1(_04985_),
    .A2(_05004_),
    .B(_05009_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10505_ (.I(_03775_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10506_ (.I(_04850_),
    .Z(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10507_ (.A1(_01517_),
    .A2(_04245_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10508_ (.A1(_03613_),
    .A2(_01617_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10509_ (.A1(_05012_),
    .A2(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10510_ (.A1(_01626_),
    .A2(_03630_),
    .B1(_03633_),
    .B2(_01604_),
    .C1(_05014_),
    .C2(_04770_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10511_ (.A1(_01617_),
    .A2(_04779_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10512_ (.A1(_01328_),
    .A2(_04954_),
    .B1(_04781_),
    .B2(_01179_),
    .C(_05016_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10513_ (.A1(_02949_),
    .A2(_01170_),
    .A3(_04773_),
    .B1(_04849_),
    .B2(_04850_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10514_ (.A1(_05011_),
    .A2(_05015_),
    .B1(_05017_),
    .B2(_05018_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10515_ (.A1(_04166_),
    .A2(_04922_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10516_ (.A1(_04963_),
    .A2(_05019_),
    .B(_05020_),
    .C(_04921_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10517_ (.A1(_02646_),
    .A2(_04811_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10518_ (.A1(_02639_),
    .A2(_01326_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10519_ (.A1(_01325_),
    .A2(_04935_),
    .B(_05023_),
    .C(_05022_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10520_ (.A1(_01618_),
    .A2(_05022_),
    .B(_05024_),
    .C(_04810_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10521_ (.A1(_01328_),
    .A2(_04940_),
    .B(_04920_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10522_ (.A1(_04940_),
    .A2(_05021_),
    .A3(_05025_),
    .B(_05026_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10523_ (.A1(_02341_),
    .A2(_04821_),
    .B(_04822_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10524_ (.A1(_05010_),
    .A2(_04877_),
    .B1(_05027_),
    .B2(_05028_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10525_ (.A1(_04166_),
    .A2(_04825_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10526_ (.A1(_04760_),
    .A2(_05029_),
    .B(_05030_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10527_ (.I(_05031_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10528_ (.I(_05032_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10529_ (.A1(_02949_),
    .A2(_04863_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10530_ (.A1(_02256_),
    .A2(_04862_),
    .B(_05034_),
    .C(_04867_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10531_ (.A1(_04108_),
    .A2(_04908_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10532_ (.A1(_05035_),
    .A2(_05036_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10533_ (.A1(\as2650.regs[5][5] ),
    .A2(_04873_),
    .B1(_05037_),
    .B2(_04871_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10534_ (.A1(_04985_),
    .A2(_05033_),
    .B(_05038_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10535_ (.A1(_01322_),
    .A2(_04954_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10536_ (.A1(_01626_),
    .A2(_04954_),
    .B(_04842_),
    .C(_05039_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10537_ (.A1(_01263_),
    .A2(_03619_),
    .A3(_03620_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10538_ (.A1(_04498_),
    .A2(_05041_),
    .B1(_04957_),
    .B2(net217),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10539_ (.A1(_01312_),
    .A2(_05012_),
    .Z(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10540_ (.A1(_04236_),
    .A2(_03630_),
    .B1(_03632_),
    .B2(_01617_),
    .C1(_05043_),
    .C2(_04770_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10541_ (.A1(_04850_),
    .A2(_05044_),
    .B(_04802_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10542_ (.A1(_05040_),
    .A2(_05042_),
    .B(_05045_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10543_ (.I(_04159_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10544_ (.A1(_05047_),
    .A2(_04797_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10545_ (.A1(_05046_),
    .A2(_05048_),
    .B(_04810_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10546_ (.A1(_02640_),
    .A2(_01320_),
    .B1(_01318_),
    .B2(_04970_),
    .C(_04934_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10547_ (.A1(_01627_),
    .A2(_05022_),
    .B(_04807_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10548_ (.A1(_05050_),
    .A2(_05051_),
    .B(_04845_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10549_ (.A1(_01323_),
    .A2(_04815_),
    .B(_04818_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10550_ (.A1(_05049_),
    .A2(_05052_),
    .B(_05053_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10551_ (.A1(_02718_),
    .A2(_04898_),
    .B(_04843_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10552_ (.A1(_03780_),
    .A2(_04843_),
    .B1(_05054_),
    .B2(_05055_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10553_ (.I0(_05056_),
    .I1(_05047_),
    .S(_04825_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10554_ (.I(_05057_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10555_ (.I(_05058_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10556_ (.A1(_04106_),
    .A2(_04908_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10557_ (.A1(_02951_),
    .A2(_04911_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10558_ (.A1(_02893_),
    .A2(_04910_),
    .B(_05061_),
    .C(_04867_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10559_ (.A1(_05060_),
    .A2(_05062_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10560_ (.A1(\as2650.regs[5][6] ),
    .A2(_04873_),
    .B1(_05063_),
    .B2(_04871_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10561_ (.A1(_04985_),
    .A2(_05059_),
    .B(_05064_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10562_ (.I(_04779_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10563_ (.A1(_01311_),
    .A2(_05065_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10564_ (.A1(_03621_),
    .A2(_05065_),
    .B1(_04781_),
    .B2(_01180_),
    .C(_05066_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10565_ (.A1(_04550_),
    .A2(_05041_),
    .B1(_04957_),
    .B2(net218),
    .C(_05067_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10566_ (.A1(_03763_),
    .A2(_04245_),
    .B(_03613_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10567_ (.A1(_01638_),
    .A2(_05069_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10568_ (.A1(_04236_),
    .A2(_05069_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10569_ (.A1(_01263_),
    .A2(_05070_),
    .A3(_05071_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10570_ (.A1(_04231_),
    .A2(_05072_),
    .B(_04550_),
    .C(_04321_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10571_ (.A1(_04963_),
    .A2(_05073_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10572_ (.A1(_03699_),
    .A2(_04963_),
    .B1(_05068_),
    .B2(_05074_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10573_ (.A1(_02640_),
    .A2(_01298_),
    .B1(_01309_),
    .B2(_04970_),
    .C(_04891_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10574_ (.A1(_01638_),
    .A2(_04891_),
    .B(_05076_),
    .C(_04921_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10575_ (.A1(_04921_),
    .A2(_05075_),
    .B(_05077_),
    .C(_04898_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10576_ (.A1(_02572_),
    .A2(_04299_),
    .B(_05078_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10577_ (.A1(_03772_),
    .A2(_04843_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10578_ (.A1(_04875_),
    .A2(_05080_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10579_ (.A1(_03700_),
    .A2(_04919_),
    .B1(_05079_),
    .B2(_05081_),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10580_ (.I(_05082_),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10581_ (.A1(_04104_),
    .A2(_04858_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10582_ (.A1(_02954_),
    .A2(_04911_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10583_ (.A1(_02924_),
    .A2(_04910_),
    .B(_05085_),
    .C(_04867_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10584_ (.A1(_05084_),
    .A2(_05086_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10585_ (.A1(\as2650.regs[5][7] ),
    .A2(_04873_),
    .B1(_05087_),
    .B2(_04871_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10586_ (.A1(_04985_),
    .A2(_05083_),
    .B(_05088_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10587_ (.A1(_04714_),
    .A2(_04629_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10588_ (.I(_05089_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10589_ (.I(_05090_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10590_ (.I(_05089_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10591_ (.I(_05092_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10592_ (.A1(\as2650.stack[2][0] ),
    .A2(_05093_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10593_ (.A1(_04713_),
    .A2(_05091_),
    .B(_05094_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10594_ (.A1(\as2650.stack[2][1] ),
    .A2(_05093_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10595_ (.A1(_04721_),
    .A2(_05091_),
    .B(_05095_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10596_ (.A1(\as2650.stack[2][2] ),
    .A2(_05093_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10597_ (.A1(_04723_),
    .A2(_05091_),
    .B(_05096_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10598_ (.A1(\as2650.stack[2][3] ),
    .A2(_05093_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10599_ (.A1(_04725_),
    .A2(_05091_),
    .B(_05097_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10600_ (.I(_05090_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10601_ (.I(_05092_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10602_ (.A1(\as2650.stack[2][4] ),
    .A2(_05099_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10603_ (.A1(_04727_),
    .A2(_05098_),
    .B(_05100_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10604_ (.A1(\as2650.stack[2][5] ),
    .A2(_05099_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10605_ (.A1(_04731_),
    .A2(_05098_),
    .B(_05101_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10606_ (.A1(\as2650.stack[2][6] ),
    .A2(_05099_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10607_ (.A1(_04733_),
    .A2(_05098_),
    .B(_05102_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10608_ (.A1(\as2650.stack[2][7] ),
    .A2(_05099_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10609_ (.A1(_04735_),
    .A2(_05098_),
    .B(_05103_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10610_ (.I(_05090_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10611_ (.I(_05092_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10612_ (.A1(\as2650.stack[2][8] ),
    .A2(_05105_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10613_ (.A1(_04737_),
    .A2(_05104_),
    .B(_05106_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10614_ (.A1(\as2650.stack[2][9] ),
    .A2(_05105_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10615_ (.A1(_04741_),
    .A2(_05104_),
    .B(_05107_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10616_ (.A1(\as2650.stack[2][10] ),
    .A2(_05105_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10617_ (.A1(_04743_),
    .A2(_05104_),
    .B(_05108_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10618_ (.A1(\as2650.stack[2][11] ),
    .A2(_05105_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10619_ (.A1(_04745_),
    .A2(_05104_),
    .B(_05109_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10620_ (.I(_05090_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10621_ (.I(_05092_),
    .Z(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10622_ (.A1(\as2650.stack[2][12] ),
    .A2(_05111_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10623_ (.A1(_04747_),
    .A2(_05110_),
    .B(_05112_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10624_ (.A1(\as2650.stack[2][13] ),
    .A2(_05111_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10625_ (.A1(_04751_),
    .A2(_05110_),
    .B(_05113_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10626_ (.A1(\as2650.stack[2][14] ),
    .A2(_05111_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10627_ (.A1(_04753_),
    .A2(_05110_),
    .B(_05114_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10628_ (.A1(\as2650.stack[2][15] ),
    .A2(_05111_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10629_ (.A1(_04755_),
    .A2(_05110_),
    .B(_05115_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10630_ (.A1(_04714_),
    .A2(_04502_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10631_ (.I(_05116_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10632_ (.I(_05117_),
    .Z(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10633_ (.I(_05116_),
    .Z(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10634_ (.I(_05119_),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10635_ (.A1(\as2650.stack[1][0] ),
    .A2(_05120_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10636_ (.A1(_04713_),
    .A2(_05118_),
    .B(_05121_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10637_ (.A1(\as2650.stack[1][1] ),
    .A2(_05120_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10638_ (.A1(_04721_),
    .A2(_05118_),
    .B(_05122_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10639_ (.A1(\as2650.stack[1][2] ),
    .A2(_05120_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10640_ (.A1(_04723_),
    .A2(_05118_),
    .B(_05123_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10641_ (.A1(\as2650.stack[1][3] ),
    .A2(_05120_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10642_ (.A1(_04725_),
    .A2(_05118_),
    .B(_05124_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10643_ (.I(_05117_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10644_ (.I(_05119_),
    .Z(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10645_ (.A1(\as2650.stack[1][4] ),
    .A2(_05126_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10646_ (.A1(_04727_),
    .A2(_05125_),
    .B(_05127_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10647_ (.A1(\as2650.stack[1][5] ),
    .A2(_05126_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10648_ (.A1(_04731_),
    .A2(_05125_),
    .B(_05128_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10649_ (.A1(\as2650.stack[1][6] ),
    .A2(_05126_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10650_ (.A1(_04733_),
    .A2(_05125_),
    .B(_05129_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(\as2650.stack[1][7] ),
    .A2(_05126_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10652_ (.A1(_04735_),
    .A2(_05125_),
    .B(_05130_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10653_ (.I(_05117_),
    .Z(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10654_ (.I(_05119_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10655_ (.A1(\as2650.stack[1][8] ),
    .A2(_05132_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10656_ (.A1(_04737_),
    .A2(_05131_),
    .B(_05133_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10657_ (.A1(\as2650.stack[1][9] ),
    .A2(_05132_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10658_ (.A1(_04741_),
    .A2(_05131_),
    .B(_05134_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10659_ (.A1(\as2650.stack[1][10] ),
    .A2(_05132_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10660_ (.A1(_04743_),
    .A2(_05131_),
    .B(_05135_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10661_ (.A1(\as2650.stack[1][11] ),
    .A2(_05132_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10662_ (.A1(_04745_),
    .A2(_05131_),
    .B(_05136_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10663_ (.I(_05117_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10664_ (.I(_05119_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10665_ (.A1(\as2650.stack[1][12] ),
    .A2(_05138_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10666_ (.A1(_04747_),
    .A2(_05137_),
    .B(_05139_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10667_ (.A1(\as2650.stack[1][13] ),
    .A2(_05138_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10668_ (.A1(_04751_),
    .A2(_05137_),
    .B(_05140_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10669_ (.A1(\as2650.stack[1][14] ),
    .A2(_05138_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10670_ (.A1(_04753_),
    .A2(_05137_),
    .B(_05141_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10671_ (.A1(\as2650.stack[1][15] ),
    .A2(_05138_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10672_ (.A1(_04755_),
    .A2(_05137_),
    .B(_05142_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10673_ (.A1(_01863_),
    .A2(_01871_),
    .A3(_04685_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10674_ (.I(_05143_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10675_ (.I(_05144_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10676_ (.I(_05143_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10677_ (.I(_05146_),
    .Z(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10678_ (.A1(\as2650.stack[15][0] ),
    .A2(_05147_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10679_ (.A1(_04713_),
    .A2(_05145_),
    .B(_05148_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10680_ (.A1(\as2650.stack[15][1] ),
    .A2(_05147_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10681_ (.A1(_04721_),
    .A2(_05145_),
    .B(_05149_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10682_ (.A1(\as2650.stack[15][2] ),
    .A2(_05147_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10683_ (.A1(_04723_),
    .A2(_05145_),
    .B(_05150_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10684_ (.A1(\as2650.stack[15][3] ),
    .A2(_05147_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10685_ (.A1(_04725_),
    .A2(_05145_),
    .B(_05151_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10686_ (.I(_05144_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10687_ (.I(_05146_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10688_ (.A1(\as2650.stack[15][4] ),
    .A2(_05153_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10689_ (.A1(_04727_),
    .A2(_05152_),
    .B(_05154_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10690_ (.A1(\as2650.stack[15][5] ),
    .A2(_05153_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10691_ (.A1(_04731_),
    .A2(_05152_),
    .B(_05155_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10692_ (.A1(\as2650.stack[15][6] ),
    .A2(_05153_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10693_ (.A1(_04733_),
    .A2(_05152_),
    .B(_05156_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10694_ (.A1(\as2650.stack[15][7] ),
    .A2(_05153_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10695_ (.A1(_04735_),
    .A2(_05152_),
    .B(_05157_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10696_ (.I(_05144_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10697_ (.I(_05146_),
    .Z(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10698_ (.A1(\as2650.stack[15][8] ),
    .A2(_05159_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10699_ (.A1(_04737_),
    .A2(_05158_),
    .B(_05160_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10700_ (.A1(\as2650.stack[15][9] ),
    .A2(_05159_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10701_ (.A1(_04741_),
    .A2(_05158_),
    .B(_05161_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10702_ (.A1(\as2650.stack[15][10] ),
    .A2(_05159_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10703_ (.A1(_04743_),
    .A2(_05158_),
    .B(_05162_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10704_ (.A1(\as2650.stack[15][11] ),
    .A2(_05159_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10705_ (.A1(_04745_),
    .A2(_05158_),
    .B(_05163_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10706_ (.I(_05144_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10707_ (.I(_05146_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10708_ (.A1(\as2650.stack[15][12] ),
    .A2(_05165_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10709_ (.A1(_04747_),
    .A2(_05164_),
    .B(_05166_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10710_ (.A1(\as2650.stack[15][13] ),
    .A2(_05165_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10711_ (.A1(_04751_),
    .A2(_05164_),
    .B(_05167_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10712_ (.A1(\as2650.stack[15][14] ),
    .A2(_05165_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10713_ (.A1(_04753_),
    .A2(_05164_),
    .B(_05168_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10714_ (.A1(\as2650.stack[15][15] ),
    .A2(_05165_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10715_ (.A1(_04755_),
    .A2(_05164_),
    .B(_05169_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10716_ (.A1(_01803_),
    .A2(_04839_),
    .A3(_04854_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10717_ (.A1(_04837_),
    .A2(_05170_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10718_ (.I(_05171_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10719_ (.A1(_01803_),
    .A2(_04837_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10720_ (.I(_05173_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10721_ (.A1(_02572_),
    .A2(_05170_),
    .A3(_05173_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10722_ (.I(_05175_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10723_ (.A1(_04869_),
    .A2(_05174_),
    .B1(_05176_),
    .B2(\as2650.regs[1][0] ),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10724_ (.A1(_04829_),
    .A2(_05172_),
    .B(_05177_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10725_ (.A1(_04915_),
    .A2(_05174_),
    .B1(_05176_),
    .B2(\as2650.regs[1][1] ),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10726_ (.A1(_04905_),
    .A2(_05172_),
    .B(_05178_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10727_ (.A1(_04951_),
    .A2(_05174_),
    .B1(_05176_),
    .B2(\as2650.regs[1][2] ),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10728_ (.A1(_04946_),
    .A2(_05172_),
    .B(_05179_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10729_ (.A1(_04983_),
    .A2(_05174_),
    .B1(_05176_),
    .B2(\as2650.regs[1][3] ),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10730_ (.A1(_04980_),
    .A2(_05172_),
    .B(_05180_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10731_ (.I(_05171_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10732_ (.I(_05173_),
    .Z(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10733_ (.I(_05175_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10734_ (.A1(_05008_),
    .A2(_05182_),
    .B1(_05183_),
    .B2(\as2650.regs[1][4] ),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10735_ (.A1(_05004_),
    .A2(_05181_),
    .B(_05184_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10736_ (.A1(_05037_),
    .A2(_05182_),
    .B1(_05183_),
    .B2(\as2650.regs[1][5] ),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10737_ (.A1(_05033_),
    .A2(_05181_),
    .B(_05185_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10738_ (.A1(_05063_),
    .A2(_05182_),
    .B1(_05183_),
    .B2(\as2650.regs[1][6] ),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10739_ (.A1(_05059_),
    .A2(_05181_),
    .B(_05186_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10740_ (.A1(_05087_),
    .A2(_05182_),
    .B1(_05183_),
    .B2(\as2650.regs[1][7] ),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10741_ (.A1(_05083_),
    .A2(_05181_),
    .B(_05187_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10742_ (.I(_04839_),
    .Z(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _10743_ (.A1(_04852_),
    .A2(_01265_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10744_ (.A1(_04539_),
    .A2(_05188_),
    .A3(_05189_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10745_ (.I(_05190_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10746_ (.I(_01442_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10747_ (.A1(_05192_),
    .A2(_05190_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10748_ (.I(_05193_),
    .Z(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10749_ (.I(\as2650.regs[2][0] ),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10750_ (.A1(_04829_),
    .A2(_05191_),
    .B1(_05194_),
    .B2(_05195_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10751_ (.I(\as2650.regs[2][1] ),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10752_ (.A1(_04905_),
    .A2(_05191_),
    .B1(_05194_),
    .B2(_05196_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10753_ (.I(\as2650.regs[2][2] ),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10754_ (.A1(_04946_),
    .A2(_05191_),
    .B1(_05194_),
    .B2(_05197_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10755_ (.I(\as2650.regs[2][3] ),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10756_ (.A1(_04980_),
    .A2(_05191_),
    .B1(_05194_),
    .B2(_05198_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10757_ (.I(_05190_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10758_ (.I(_05193_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10759_ (.A1(_05004_),
    .A2(_05199_),
    .B1(_05200_),
    .B2(_00825_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10760_ (.A1(_05033_),
    .A2(_05199_),
    .B1(_05200_),
    .B2(_00844_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10761_ (.A1(_05059_),
    .A2(_05199_),
    .B1(_05200_),
    .B2(_00882_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10762_ (.A1(_05083_),
    .A2(_05199_),
    .B1(_05200_),
    .B2(_00703_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10763_ (.I(_04493_),
    .Z(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10764_ (.A1(_04381_),
    .A2(_04267_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10765_ (.A1(_04657_),
    .A2(_05202_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10766_ (.I(_05203_),
    .Z(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10767_ (.I(_05204_),
    .Z(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10768_ (.I(_05203_),
    .Z(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10769_ (.I(_05206_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10770_ (.A1(\as2650.stack[8][0] ),
    .A2(_05207_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10771_ (.A1(_05201_),
    .A2(_05205_),
    .B(_05208_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10772_ (.I(_04517_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(\as2650.stack[8][1] ),
    .A2(_05207_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10774_ (.A1(_05209_),
    .A2(_05205_),
    .B(_05210_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10775_ (.I(_04525_),
    .Z(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10776_ (.A1(\as2650.stack[8][2] ),
    .A2(_05207_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10777_ (.A1(_05211_),
    .A2(_05205_),
    .B(_05212_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10778_ (.I(_04533_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(\as2650.stack[8][3] ),
    .A2(_05207_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10780_ (.A1(_05213_),
    .A2(_05205_),
    .B(_05214_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10781_ (.I(_04543_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10782_ (.I(_05204_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10783_ (.I(_05206_),
    .Z(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10784_ (.A1(\as2650.stack[8][4] ),
    .A2(_05217_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10785_ (.A1(_05215_),
    .A2(_05216_),
    .B(_05218_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10786_ (.I(_04556_),
    .Z(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10787_ (.A1(\as2650.stack[8][5] ),
    .A2(_05217_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10788_ (.A1(_05219_),
    .A2(_05216_),
    .B(_05220_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10789_ (.I(_04563_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10790_ (.A1(\as2650.stack[8][6] ),
    .A2(_05217_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10791_ (.A1(_05221_),
    .A2(_05216_),
    .B(_05222_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10792_ (.I(_04570_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10793_ (.A1(\as2650.stack[8][7] ),
    .A2(_05217_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10794_ (.A1(_05223_),
    .A2(_05216_),
    .B(_05224_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10795_ (.I(_04578_),
    .Z(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10796_ (.I(_05204_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10797_ (.I(_05206_),
    .Z(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10798_ (.A1(\as2650.stack[8][8] ),
    .A2(_05227_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10799_ (.A1(_05225_),
    .A2(_05226_),
    .B(_05228_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10800_ (.I(_04586_),
    .Z(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10801_ (.A1(\as2650.stack[8][9] ),
    .A2(_05227_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10802_ (.A1(_05229_),
    .A2(_05226_),
    .B(_05230_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10803_ (.I(_04594_),
    .Z(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10804_ (.A1(\as2650.stack[8][10] ),
    .A2(_05227_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10805_ (.A1(_05231_),
    .A2(_05226_),
    .B(_05232_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10806_ (.I(_04600_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10807_ (.A1(\as2650.stack[8][11] ),
    .A2(_05227_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10808_ (.A1(_05233_),
    .A2(_05226_),
    .B(_05234_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10809_ (.I(_04607_),
    .Z(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10810_ (.I(_05204_),
    .Z(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10811_ (.I(_05206_),
    .Z(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10812_ (.A1(\as2650.stack[8][12] ),
    .A2(_05237_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10813_ (.A1(_05235_),
    .A2(_05236_),
    .B(_05238_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10814_ (.I(_04615_),
    .Z(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10815_ (.A1(\as2650.stack[8][13] ),
    .A2(_05237_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10816_ (.A1(_05239_),
    .A2(_05236_),
    .B(_05240_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10817_ (.I(_04621_),
    .Z(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10818_ (.A1(\as2650.stack[8][14] ),
    .A2(_05237_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10819_ (.A1(_05241_),
    .A2(_05236_),
    .B(_05242_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10820_ (.I(_04626_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10821_ (.A1(\as2650.stack[8][15] ),
    .A2(_05237_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10822_ (.A1(_05243_),
    .A2(_05236_),
    .B(_05244_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10823_ (.A1(_04539_),
    .A2(_05188_),
    .A3(_04853_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10824_ (.I(_05245_),
    .Z(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10825_ (.A1(_05192_),
    .A2(_05245_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10826_ (.I(_05247_),
    .Z(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10827_ (.A1(_04829_),
    .A2(_05246_),
    .B1(_05248_),
    .B2(_00737_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10828_ (.A1(_04905_),
    .A2(_05246_),
    .B1(_05248_),
    .B2(_00754_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10829_ (.A1(_04946_),
    .A2(_05246_),
    .B1(_05248_),
    .B2(_00779_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10830_ (.A1(_04980_),
    .A2(_05246_),
    .B1(_05248_),
    .B2(_00801_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10831_ (.I(_05245_),
    .Z(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10832_ (.I(_05247_),
    .Z(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10833_ (.A1(_05004_),
    .A2(_05249_),
    .B1(_05250_),
    .B2(_00829_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10834_ (.A1(_05033_),
    .A2(_05249_),
    .B1(_05250_),
    .B2(_00847_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10835_ (.A1(_05059_),
    .A2(_05249_),
    .B1(_05250_),
    .B2(_00885_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10836_ (.A1(_05083_),
    .A2(_05249_),
    .B1(_05250_),
    .B2(_00708_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10837_ (.A1(_00148_),
    .A2(_01542_),
    .A3(_01545_),
    .Z(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10838_ (.I(_05251_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10839_ (.A1(_03735_),
    .A2(_05188_),
    .A3(_05189_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10840_ (.I(_05252_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10841_ (.A1(_05192_),
    .A2(_05252_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10842_ (.I(_05254_),
    .Z(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10843_ (.I(\as2650.regs[6][0] ),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10844_ (.A1(_04828_),
    .A2(_05253_),
    .B1(_05255_),
    .B2(_05256_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10845_ (.I(\as2650.regs[6][1] ),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10846_ (.A1(_04904_),
    .A2(_05253_),
    .B1(_05255_),
    .B2(_05257_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10847_ (.I(\as2650.regs[6][2] ),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10848_ (.A1(_04945_),
    .A2(_05253_),
    .B1(_05255_),
    .B2(_05258_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10849_ (.I(_04979_),
    .Z(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10850_ (.I(\as2650.regs[6][3] ),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10851_ (.A1(_05259_),
    .A2(_05253_),
    .B1(_05255_),
    .B2(_05260_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10852_ (.I(_05252_),
    .Z(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10853_ (.I(_05254_),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10854_ (.I(\as2650.regs[6][4] ),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10855_ (.A1(_05003_),
    .A2(_05261_),
    .B1(_05262_),
    .B2(_05263_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10856_ (.I(\as2650.regs[6][5] ),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10857_ (.A1(_05032_),
    .A2(_05261_),
    .B1(_05262_),
    .B2(_05264_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10858_ (.I(\as2650.regs[6][6] ),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10859_ (.A1(_05058_),
    .A2(_05261_),
    .B1(_05262_),
    .B2(_05265_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10860_ (.I(_05082_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10861_ (.I(\as2650.regs[6][7] ),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10862_ (.A1(_05266_),
    .A2(_05261_),
    .B1(_05262_),
    .B2(_05267_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10863_ (.A1(_02876_),
    .A2(_04714_),
    .A3(_04500_),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10864_ (.I(_05268_),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10865_ (.I(_05269_),
    .Z(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10866_ (.I(_05268_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10867_ (.I(_05271_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10868_ (.A1(\as2650.stack[0][0] ),
    .A2(_05272_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10869_ (.A1(_05201_),
    .A2(_05270_),
    .B(_05273_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10870_ (.A1(\as2650.stack[0][1] ),
    .A2(_05272_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10871_ (.A1(_05209_),
    .A2(_05270_),
    .B(_05274_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10872_ (.A1(\as2650.stack[0][2] ),
    .A2(_05272_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10873_ (.A1(_05211_),
    .A2(_05270_),
    .B(_05275_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10874_ (.A1(\as2650.stack[0][3] ),
    .A2(_05272_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10875_ (.A1(_05213_),
    .A2(_05270_),
    .B(_05276_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10876_ (.I(_05269_),
    .Z(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10877_ (.I(_05271_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10878_ (.A1(\as2650.stack[0][4] ),
    .A2(_05278_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10879_ (.A1(_05215_),
    .A2(_05277_),
    .B(_05279_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10880_ (.A1(\as2650.stack[0][5] ),
    .A2(_05278_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10881_ (.A1(_05219_),
    .A2(_05277_),
    .B(_05280_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10882_ (.A1(\as2650.stack[0][6] ),
    .A2(_05278_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10883_ (.A1(_05221_),
    .A2(_05277_),
    .B(_05281_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10884_ (.A1(\as2650.stack[0][7] ),
    .A2(_05278_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10885_ (.A1(_05223_),
    .A2(_05277_),
    .B(_05282_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10886_ (.I(_05269_),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10887_ (.I(_05271_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10888_ (.A1(\as2650.stack[0][8] ),
    .A2(_05284_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10889_ (.A1(_05225_),
    .A2(_05283_),
    .B(_05285_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10890_ (.A1(\as2650.stack[0][9] ),
    .A2(_05284_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10891_ (.A1(_05229_),
    .A2(_05283_),
    .B(_05286_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10892_ (.A1(\as2650.stack[0][10] ),
    .A2(_05284_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10893_ (.A1(_05231_),
    .A2(_05283_),
    .B(_05287_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10894_ (.A1(\as2650.stack[0][11] ),
    .A2(_05284_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10895_ (.A1(_05233_),
    .A2(_05283_),
    .B(_05288_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10896_ (.I(_05269_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10897_ (.I(_05271_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10898_ (.A1(\as2650.stack[0][12] ),
    .A2(_05290_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10899_ (.A1(_05235_),
    .A2(_05289_),
    .B(_05291_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10900_ (.A1(\as2650.stack[0][13] ),
    .A2(_05290_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10901_ (.A1(_05239_),
    .A2(_05289_),
    .B(_05292_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10902_ (.A1(\as2650.stack[0][14] ),
    .A2(_05290_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10903_ (.A1(_05241_),
    .A2(_05289_),
    .B(_05293_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10904_ (.A1(\as2650.stack[0][15] ),
    .A2(_05290_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10905_ (.A1(_05243_),
    .A2(_05289_),
    .B(_05294_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10906_ (.A1(_04685_),
    .A2(_05202_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10907_ (.I(_05295_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10908_ (.I(_05296_),
    .Z(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10909_ (.I(_05295_),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10910_ (.I(_05298_),
    .Z(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10911_ (.A1(\as2650.stack[11][0] ),
    .A2(_05299_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10912_ (.A1(_05201_),
    .A2(_05297_),
    .B(_05300_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10913_ (.A1(\as2650.stack[11][1] ),
    .A2(_05299_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10914_ (.A1(_05209_),
    .A2(_05297_),
    .B(_05301_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10915_ (.A1(\as2650.stack[11][2] ),
    .A2(_05299_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10916_ (.A1(_05211_),
    .A2(_05297_),
    .B(_05302_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10917_ (.A1(\as2650.stack[11][3] ),
    .A2(_05299_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10918_ (.A1(_05213_),
    .A2(_05297_),
    .B(_05303_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10919_ (.I(_05296_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10920_ (.I(_05298_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10921_ (.A1(\as2650.stack[11][4] ),
    .A2(_05305_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10922_ (.A1(_05215_),
    .A2(_05304_),
    .B(_05306_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10923_ (.A1(\as2650.stack[11][5] ),
    .A2(_05305_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10924_ (.A1(_05219_),
    .A2(_05304_),
    .B(_05307_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10925_ (.A1(\as2650.stack[11][6] ),
    .A2(_05305_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10926_ (.A1(_05221_),
    .A2(_05304_),
    .B(_05308_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10927_ (.A1(\as2650.stack[11][7] ),
    .A2(_05305_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10928_ (.A1(_05223_),
    .A2(_05304_),
    .B(_05309_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10929_ (.I(_05296_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10930_ (.I(_05298_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10931_ (.A1(\as2650.stack[11][8] ),
    .A2(_05311_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10932_ (.A1(_05225_),
    .A2(_05310_),
    .B(_05312_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10933_ (.A1(\as2650.stack[11][9] ),
    .A2(_05311_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10934_ (.A1(_05229_),
    .A2(_05310_),
    .B(_05313_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10935_ (.A1(\as2650.stack[11][10] ),
    .A2(_05311_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10936_ (.A1(_05231_),
    .A2(_05310_),
    .B(_05314_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10937_ (.A1(\as2650.stack[11][11] ),
    .A2(_05311_),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10938_ (.A1(_05233_),
    .A2(_05310_),
    .B(_05315_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10939_ (.I(_05296_),
    .Z(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10940_ (.I(_05298_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10941_ (.A1(\as2650.stack[11][12] ),
    .A2(_05317_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10942_ (.A1(_05235_),
    .A2(_05316_),
    .B(_05318_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10943_ (.A1(\as2650.stack[11][13] ),
    .A2(_05317_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10944_ (.A1(_05239_),
    .A2(_05316_),
    .B(_05319_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10945_ (.A1(\as2650.stack[11][14] ),
    .A2(_05317_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10946_ (.A1(_05241_),
    .A2(_05316_),
    .B(_05320_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10947_ (.A1(\as2650.stack[11][15] ),
    .A2(_05317_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10948_ (.A1(_05243_),
    .A2(_05316_),
    .B(_05321_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10949_ (.I(_01802_),
    .Z(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10950_ (.A1(_02270_),
    .A2(_02932_),
    .A3(_04431_),
    .A4(_04780_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10951_ (.A1(_01180_),
    .A2(_05323_),
    .B(_04832_),
    .C(_04830_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10952_ (.A1(_03626_),
    .A2(_04484_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10953_ (.A1(_04311_),
    .A2(_04550_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10954_ (.A1(_01537_),
    .A2(_04771_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10955_ (.I(_05327_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10956_ (.A1(_05324_),
    .A2(_05325_),
    .A3(_05326_),
    .A4(_05328_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10957_ (.A1(_05322_),
    .A2(_05329_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10958_ (.I(_05330_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10959_ (.A1(_03806_),
    .A2(_05011_),
    .ZN(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10960_ (.I(_05332_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10961_ (.I(_05333_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10962_ (.I(_05328_),
    .Z(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10963_ (.I(_04833_),
    .Z(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10964_ (.I(_05327_),
    .Z(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10965_ (.A1(_03000_),
    .A2(_05336_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10966_ (.A1(_02956_),
    .A2(_05336_),
    .B(_05337_),
    .C(_05338_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10967_ (.I(_04948_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10968_ (.A1(\as2650.chirpchar[0] ),
    .A2(_05335_),
    .B(_05339_),
    .C(_05340_),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10969_ (.A1(net219),
    .A2(net188),
    .A3(_04858_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10970_ (.A1(_03638_),
    .A2(_05011_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10971_ (.I(_05343_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10972_ (.I(_05344_),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10973_ (.A1(_05341_),
    .A2(_05342_),
    .B(_05345_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10974_ (.I(_05325_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10975_ (.A1(_04199_),
    .A2(_05347_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10976_ (.I(_05332_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10977_ (.A1(_04273_),
    .A2(_05349_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10978_ (.A1(_05334_),
    .A2(_05346_),
    .A3(_05348_),
    .B(_05350_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10979_ (.A1(_01629_),
    .A2(_04758_),
    .B(_05189_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10980_ (.A1(_03730_),
    .A2(_04838_),
    .A3(_05352_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10981_ (.I(_05329_),
    .Z(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10982_ (.A1(_03731_),
    .A2(_01659_),
    .A3(_05353_),
    .A4(_05354_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10983_ (.I(_05355_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10984_ (.A1(\as2650.regs[4][0] ),
    .A2(_05356_),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10985_ (.I(_05322_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10986_ (.I(_01659_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _10987_ (.A1(_00691_),
    .A2(_04838_),
    .A3(_05352_),
    .Z(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10988_ (.A1(_05358_),
    .A2(_00724_),
    .A3(_05359_),
    .B1(_04827_),
    .B2(_05360_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10989_ (.I(_05330_),
    .Z(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10990_ (.A1(_05361_),
    .A2(_05362_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10991_ (.A1(_05331_),
    .A2(_05351_),
    .B(_05357_),
    .C(_05363_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10992_ (.I(_05326_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10993_ (.I(_05325_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10994_ (.A1(_04128_),
    .A2(_04907_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10995_ (.I(_04832_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10996_ (.A1(_03063_),
    .A2(_05367_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10997_ (.A1(_00749_),
    .A2(_04834_),
    .B(_05328_),
    .C(_05368_),
    .ZN(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10998_ (.A1(\as2650.chirpchar[1] ),
    .A2(_05337_),
    .B(_05369_),
    .C(_04948_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10999_ (.A1(_04002_),
    .A2(_05366_),
    .B(_05370_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11000_ (.A1(_05365_),
    .A2(_05371_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11001_ (.A1(_04192_),
    .A2(_05347_),
    .B(_05364_),
    .C(_05372_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11002_ (.A1(_04279_),
    .A2(_05334_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11003_ (.A1(_05373_),
    .A2(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11004_ (.A1(\as2650.regs[4][1] ),
    .A2(_05356_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11005_ (.I(_05330_),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11006_ (.I(_03735_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11007_ (.I(_05360_),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11008_ (.A1(_05378_),
    .A2(_00745_),
    .A3(_02573_),
    .B1(_04903_),
    .B2(_05379_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11009_ (.A1(_05377_),
    .A2(_05380_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11010_ (.A1(_05331_),
    .A2(_05375_),
    .B(_05376_),
    .C(_05381_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _11011_ (.A1(_05324_),
    .A2(_05325_),
    .A3(_05326_),
    .A4(_05335_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11012_ (.A1(_03732_),
    .A2(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11013_ (.A1(_04918_),
    .A2(_04919_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11014_ (.A1(_04919_),
    .A2(_04943_),
    .B(_05384_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11015_ (.A1(_05359_),
    .A2(_05353_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11016_ (.A1(_05385_),
    .A2(_05353_),
    .B1(_05386_),
    .B2(_00769_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11017_ (.I(_05355_),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11018_ (.A1(\as2650.regs[4][2] ),
    .A2(_05388_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11019_ (.I(_05327_),
    .Z(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11020_ (.A1(_03105_),
    .A2(_04833_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11021_ (.A1(_00772_),
    .A2(_05367_),
    .B(_05327_),
    .C(_05391_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11022_ (.A1(\as2650.chirpchar[2] ),
    .A2(_05390_),
    .B(_05392_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11023_ (.A1(_04866_),
    .A2(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11024_ (.A1(_04127_),
    .A2(_05340_),
    .B(_05365_),
    .C(_05394_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11025_ (.A1(_04183_),
    .A2(_05347_),
    .B(_05364_),
    .C(_05395_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11026_ (.A1(_04265_),
    .A2(_05349_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11027_ (.A1(_05396_),
    .A2(_05397_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11028_ (.A1(_05362_),
    .A2(_05398_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11029_ (.A1(_05383_),
    .A2(_05387_),
    .B(_05389_),
    .C(_05399_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11030_ (.A1(_04539_),
    .A2(\as2650.regs[0][3] ),
    .A3(_02138_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11031_ (.A1(_05259_),
    .A2(_05379_),
    .B(_05400_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11032_ (.A1(_05377_),
    .A2(_05401_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11033_ (.A1(_03142_),
    .A2(_04834_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11034_ (.A1(_00796_),
    .A2(_05336_),
    .B(_05390_),
    .C(_05403_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11035_ (.A1(\as2650.chirpchar[3] ),
    .A2(_05335_),
    .B(_05404_),
    .C(_05340_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11036_ (.A1(_04125_),
    .A2(_04949_),
    .B(_05365_),
    .C(_05405_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11037_ (.A1(_04175_),
    .A2(_05345_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11038_ (.A1(_05364_),
    .A2(_05406_),
    .A3(_05407_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11039_ (.A1(_04269_),
    .A2(_05349_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11040_ (.A1(_05408_),
    .A2(_05409_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11041_ (.A1(\as2650.regs[4][3] ),
    .A2(_05356_),
    .B1(_05410_),
    .B2(_05383_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11042_ (.A1(_05402_),
    .A2(_05411_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11043_ (.A1(_03186_),
    .A2(_05367_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11044_ (.A1(_00822_),
    .A2(_04834_),
    .B(_05390_),
    .C(_05412_),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11045_ (.A1(\as2650.chirpchar[4] ),
    .A2(_05335_),
    .B(_05413_),
    .C(_04866_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11046_ (.A1(_04124_),
    .A2(_04949_),
    .B(_05365_),
    .C(_05414_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11047_ (.A1(_03754_),
    .A2(_05347_),
    .B(_05415_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11048_ (.I0(_04281_),
    .I1(_05416_),
    .S(_05364_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11049_ (.A1(\as2650.regs[4][4] ),
    .A2(_05388_),
    .ZN(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11050_ (.A1(_05378_),
    .A2(_00814_),
    .A3(_02573_),
    .B1(_05002_),
    .B2(_05379_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11051_ (.A1(_05377_),
    .A2(_05419_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11052_ (.A1(_05331_),
    .A2(_05417_),
    .B(_05418_),
    .C(_05420_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11053_ (.A1(_04275_),
    .A2(_04276_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11054_ (.A1(_03223_),
    .A2(_04833_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11055_ (.A1(_02967_),
    .A2(_05367_),
    .B(_05328_),
    .C(_05422_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11056_ (.A1(\as2650.chirpchar[5] ),
    .A2(_05337_),
    .B(_05423_),
    .C(_04948_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11057_ (.A1(_04122_),
    .A2(_05340_),
    .B(_05424_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11058_ (.A1(_05344_),
    .A2(_05425_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11059_ (.A1(_04166_),
    .A2(_05345_),
    .B(_05333_),
    .C(_05426_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11060_ (.A1(_05421_),
    .A2(_05334_),
    .B(_05427_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11061_ (.A1(\as2650.regs[4][5] ),
    .A2(_05388_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11062_ (.A1(_05358_),
    .A2(_00852_),
    .A3(_05359_),
    .B1(_05031_),
    .B2(_05360_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11063_ (.A1(_05362_),
    .A2(_05430_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11064_ (.A1(_05331_),
    .A2(_05428_),
    .B(_05429_),
    .C(_05431_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11065_ (.A1(_02969_),
    .A2(_04860_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11066_ (.A1(_03257_),
    .A2(_04860_),
    .B(_05432_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11067_ (.A1(\as2650.chirpchar[6] ),
    .A2(_05390_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11068_ (.A1(_05337_),
    .A2(_05433_),
    .B(_05434_),
    .C(_04907_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11069_ (.A1(_04120_),
    .A2(_04858_),
    .B(_05344_),
    .C(_05435_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11070_ (.A1(_05047_),
    .A2(_05345_),
    .B(_05333_),
    .C(_05436_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11071_ (.A1(_04270_),
    .A2(_05334_),
    .B(_05437_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11072_ (.A1(_05358_),
    .A2(_00872_),
    .A3(_05359_),
    .B1(_05057_),
    .B2(_05360_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11073_ (.A1(_05362_),
    .A2(_05439_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11074_ (.A1(\as2650.regs[4][6] ),
    .A2(_05356_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11075_ (.A1(_05377_),
    .A2(_05438_),
    .B(_05440_),
    .C(_05441_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11076_ (.I(_03296_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11077_ (.A1(_05442_),
    .A2(_04831_),
    .B(_04139_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11078_ (.A1(net194),
    .A2(_05336_),
    .B1(_05443_),
    .B2(_05011_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11079_ (.A1(_04119_),
    .A2(_04907_),
    .B(_05343_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11080_ (.A1(_03699_),
    .A2(_05344_),
    .B1(_05444_),
    .B2(_05445_),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11081_ (.A1(_05333_),
    .A2(_05446_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11082_ (.A1(_04261_),
    .A2(_05349_),
    .B(_05382_),
    .C(_05447_),
    .ZN(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11083_ (.A1(_00692_),
    .A2(_05386_),
    .B1(_05388_),
    .B2(\as2650.regs[4][7] ),
    .C1(_05378_),
    .C2(_05448_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11084_ (.A1(_05266_),
    .A2(_05379_),
    .A3(_05354_),
    .B(_05449_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11085_ (.A1(_04629_),
    .A2(_05202_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11086_ (.I(_05450_),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11087_ (.I(_05451_),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11088_ (.I(_05450_),
    .Z(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11089_ (.I(_05453_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11090_ (.A1(\as2650.stack[10][0] ),
    .A2(_05454_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11091_ (.A1(_05201_),
    .A2(_05452_),
    .B(_05455_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11092_ (.A1(\as2650.stack[10][1] ),
    .A2(_05454_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11093_ (.A1(_05209_),
    .A2(_05452_),
    .B(_05456_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11094_ (.A1(\as2650.stack[10][2] ),
    .A2(_05454_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11095_ (.A1(_05211_),
    .A2(_05452_),
    .B(_05457_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11096_ (.A1(\as2650.stack[10][3] ),
    .A2(_05454_),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11097_ (.A1(_05213_),
    .A2(_05452_),
    .B(_05458_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11098_ (.I(_05451_),
    .Z(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11099_ (.I(_05453_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11100_ (.A1(\as2650.stack[10][4] ),
    .A2(_05460_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11101_ (.A1(_05215_),
    .A2(_05459_),
    .B(_05461_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11102_ (.A1(\as2650.stack[10][5] ),
    .A2(_05460_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11103_ (.A1(_05219_),
    .A2(_05459_),
    .B(_05462_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11104_ (.A1(\as2650.stack[10][6] ),
    .A2(_05460_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11105_ (.A1(_05221_),
    .A2(_05459_),
    .B(_05463_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11106_ (.A1(\as2650.stack[10][7] ),
    .A2(_05460_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11107_ (.A1(_05223_),
    .A2(_05459_),
    .B(_05464_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11108_ (.I(_05451_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11109_ (.I(_05453_),
    .Z(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11110_ (.A1(\as2650.stack[10][8] ),
    .A2(_05466_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11111_ (.A1(_05225_),
    .A2(_05465_),
    .B(_05467_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11112_ (.A1(\as2650.stack[10][9] ),
    .A2(_05466_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11113_ (.A1(_05229_),
    .A2(_05465_),
    .B(_05468_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11114_ (.A1(\as2650.stack[10][10] ),
    .A2(_05466_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11115_ (.A1(_05231_),
    .A2(_05465_),
    .B(_05469_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11116_ (.A1(\as2650.stack[10][11] ),
    .A2(_05466_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11117_ (.A1(_05233_),
    .A2(_05465_),
    .B(_05470_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11118_ (.I(_05451_),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11119_ (.I(_05453_),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11120_ (.A1(\as2650.stack[10][12] ),
    .A2(_05472_),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11121_ (.A1(_05235_),
    .A2(_05471_),
    .B(_05473_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11122_ (.A1(\as2650.stack[10][13] ),
    .A2(_05472_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11123_ (.A1(_05239_),
    .A2(_05471_),
    .B(_05474_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11124_ (.A1(\as2650.stack[10][14] ),
    .A2(_05472_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11125_ (.A1(_05241_),
    .A2(_05471_),
    .B(_05475_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11126_ (.A1(\as2650.stack[10][15] ),
    .A2(_05472_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11127_ (.A1(_05243_),
    .A2(_05471_),
    .B(_05476_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11128_ (.A1(_03731_),
    .A2(_05329_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11129_ (.I(_05477_),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _11130_ (.A1(_01802_),
    .A2(_04838_),
    .A3(_05352_),
    .Z(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11131_ (.I(_01550_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11132_ (.A1(_01804_),
    .A2(\as2650.regs[4][0] ),
    .A3(_05480_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11133_ (.A1(_04828_),
    .A2(_05479_),
    .B(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11134_ (.I(_05477_),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11135_ (.A1(_05482_),
    .A2(_05483_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11136_ (.A1(_01803_),
    .A2(_04839_),
    .A3(_05352_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11137_ (.A1(_05322_),
    .A2(_01659_),
    .A3(_05354_),
    .A4(_05485_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11138_ (.I(_05486_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11139_ (.A1(\as2650.regs[0][0] ),
    .A2(_05487_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11140_ (.A1(_05351_),
    .A2(_05478_),
    .B(_05484_),
    .C(_05488_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11141_ (.I(_05477_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11142_ (.I(_05479_),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11143_ (.I(_05322_),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11144_ (.A1(_05491_),
    .A2(\as2650.regs[4][1] ),
    .A3(_05480_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11145_ (.A1(_04904_),
    .A2(_05490_),
    .B(_05492_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11146_ (.A1(_05489_),
    .A2(_05493_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11147_ (.A1(\as2650.regs[0][1] ),
    .A2(_05487_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11148_ (.A1(_05375_),
    .A2(_05478_),
    .B(_05494_),
    .C(_05495_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11149_ (.A1(_05378_),
    .A2(_05382_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11150_ (.A1(_01804_),
    .A2(\as2650.regs[4][2] ),
    .A3(_01508_),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11151_ (.A1(_05385_),
    .A2(_05485_),
    .B(_05497_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11152_ (.I(_05486_),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11153_ (.A1(\as2650.regs[0][2] ),
    .A2(_05499_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11154_ (.A1(_05398_),
    .A2(_05489_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11155_ (.A1(_05496_),
    .A2(_05498_),
    .B(_05500_),
    .C(_05501_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11156_ (.A1(_05358_),
    .A2(\as2650.regs[4][3] ),
    .A3(_02138_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11157_ (.A1(_05259_),
    .A2(_05490_),
    .B(_05502_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11158_ (.A1(_05483_),
    .A2(_05503_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11159_ (.A1(_05410_),
    .A2(_05496_),
    .B1(_05499_),
    .B2(\as2650.regs[0][3] ),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11160_ (.A1(_05504_),
    .A2(_05505_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11161_ (.A1(_05491_),
    .A2(\as2650.regs[4][4] ),
    .A3(_05480_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11162_ (.A1(_05003_),
    .A2(_05479_),
    .B(_05506_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11163_ (.A1(_05489_),
    .A2(_05507_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11164_ (.A1(\as2650.regs[0][4] ),
    .A2(_05487_),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11165_ (.A1(_05417_),
    .A2(_05478_),
    .B(_05508_),
    .C(_05509_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11166_ (.A1(_05491_),
    .A2(\as2650.regs[4][5] ),
    .A3(_05480_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11167_ (.A1(_05032_),
    .A2(_05479_),
    .B(_05510_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11168_ (.A1(_05489_),
    .A2(_05511_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11169_ (.A1(\as2650.regs[0][5] ),
    .A2(_05487_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11170_ (.A1(_05428_),
    .A2(_05478_),
    .B(_05512_),
    .C(_05513_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11171_ (.A1(\as2650.regs[0][6] ),
    .A2(_05499_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11172_ (.A1(_05491_),
    .A2(\as2650.regs[4][6] ),
    .A3(_01508_),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11173_ (.A1(_05058_),
    .A2(_05490_),
    .B(_05515_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11174_ (.A1(_05483_),
    .A2(_05516_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11175_ (.A1(_05438_),
    .A2(_05483_),
    .B(_05514_),
    .C(_05517_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11176_ (.A1(_01804_),
    .A2(\as2650.regs[4][7] ),
    .A3(_02630_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11177_ (.A1(_03732_),
    .A2(_05448_),
    .B1(_05499_),
    .B2(\as2650.regs[0][7] ),
    .C(_05518_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11178_ (.A1(_05266_),
    .A2(_05354_),
    .A3(_05490_),
    .B(_05519_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11179_ (.A1(_03735_),
    .A2(_05188_),
    .A3(_04853_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11180_ (.I(_05520_),
    .Z(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11181_ (.A1(_05192_),
    .A2(_05520_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11182_ (.I(_05522_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11183_ (.I(\as2650.regs[7][0] ),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11184_ (.A1(_04828_),
    .A2(_05521_),
    .B1(_05523_),
    .B2(_05524_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11185_ (.I(\as2650.regs[7][1] ),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11186_ (.A1(_04904_),
    .A2(_05521_),
    .B1(_05523_),
    .B2(_05525_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11187_ (.I(\as2650.regs[7][2] ),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11188_ (.A1(_04945_),
    .A2(_05521_),
    .B1(_05523_),
    .B2(_05526_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11189_ (.I(\as2650.regs[7][3] ),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11190_ (.A1(_05259_),
    .A2(_05521_),
    .B1(_05523_),
    .B2(_05527_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11191_ (.I(_05520_),
    .Z(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11192_ (.I(_05522_),
    .Z(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11193_ (.I(\as2650.regs[7][4] ),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11194_ (.A1(_05003_),
    .A2(_05528_),
    .B1(_05529_),
    .B2(_05530_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11195_ (.I(\as2650.regs[7][5] ),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11196_ (.A1(_05032_),
    .A2(_05528_),
    .B1(_05529_),
    .B2(_05531_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11197_ (.I(\as2650.regs[7][6] ),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11198_ (.A1(_05058_),
    .A2(_05528_),
    .B1(_05529_),
    .B2(_05532_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11199_ (.I(\as2650.regs[7][7] ),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11200_ (.A1(_05266_),
    .A2(_05528_),
    .B1(_05529_),
    .B2(_05533_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11201_ (.I(_04493_),
    .Z(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11202_ (.A1(_01863_),
    .A2(_04495_),
    .A3(_04629_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11203_ (.I(_05535_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11204_ (.I(_05536_),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11205_ (.I(_05535_),
    .Z(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11206_ (.I(_05538_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11207_ (.A1(\as2650.stack[14][0] ),
    .A2(_05539_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11208_ (.A1(_05534_),
    .A2(_05537_),
    .B(_05540_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11209_ (.I(_04517_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11210_ (.A1(\as2650.stack[14][1] ),
    .A2(_05539_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11211_ (.A1(_05541_),
    .A2(_05537_),
    .B(_05542_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11212_ (.I(_04525_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11213_ (.A1(\as2650.stack[14][2] ),
    .A2(_05539_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11214_ (.A1(_05543_),
    .A2(_05537_),
    .B(_05544_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11215_ (.I(_04533_),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11216_ (.A1(\as2650.stack[14][3] ),
    .A2(_05539_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11217_ (.A1(_05545_),
    .A2(_05537_),
    .B(_05546_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11218_ (.I(_04543_),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11219_ (.I(_05536_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11220_ (.I(_05538_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11221_ (.A1(\as2650.stack[14][4] ),
    .A2(_05549_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11222_ (.A1(_05547_),
    .A2(_05548_),
    .B(_05550_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11223_ (.I(_04556_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11224_ (.A1(\as2650.stack[14][5] ),
    .A2(_05549_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11225_ (.A1(_05551_),
    .A2(_05548_),
    .B(_05552_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11226_ (.I(_04563_),
    .Z(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11227_ (.A1(\as2650.stack[14][6] ),
    .A2(_05549_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11228_ (.A1(_05553_),
    .A2(_05548_),
    .B(_05554_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11229_ (.I(_04570_),
    .Z(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11230_ (.A1(\as2650.stack[14][7] ),
    .A2(_05549_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11231_ (.A1(_05555_),
    .A2(_05548_),
    .B(_05556_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11232_ (.I(_04578_),
    .Z(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11233_ (.I(_05536_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11234_ (.I(_05538_),
    .Z(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11235_ (.A1(\as2650.stack[14][8] ),
    .A2(_05559_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11236_ (.A1(_05557_),
    .A2(_05558_),
    .B(_05560_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11237_ (.I(_04586_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11238_ (.A1(\as2650.stack[14][9] ),
    .A2(_05559_),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11239_ (.A1(_05561_),
    .A2(_05558_),
    .B(_05562_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11240_ (.I(_04594_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11241_ (.A1(\as2650.stack[14][10] ),
    .A2(_05559_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11242_ (.A1(_05563_),
    .A2(_05558_),
    .B(_05564_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11243_ (.I(_04600_),
    .Z(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11244_ (.A1(\as2650.stack[14][11] ),
    .A2(_05559_),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11245_ (.A1(_05565_),
    .A2(_05558_),
    .B(_05566_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11246_ (.I(_04607_),
    .Z(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11247_ (.I(_05536_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11248_ (.I(_05538_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11249_ (.A1(\as2650.stack[14][12] ),
    .A2(_05569_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11250_ (.A1(_05567_),
    .A2(_05568_),
    .B(_05570_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11251_ (.I(_04615_),
    .Z(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11252_ (.A1(\as2650.stack[14][13] ),
    .A2(_05569_),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11253_ (.A1(_05571_),
    .A2(_05568_),
    .B(_05572_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11254_ (.I(_04621_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11255_ (.A1(\as2650.stack[14][14] ),
    .A2(_05569_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11256_ (.A1(_05573_),
    .A2(_05568_),
    .B(_05574_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11257_ (.I(_04626_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11258_ (.A1(\as2650.stack[14][15] ),
    .A2(_05569_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11259_ (.A1(_05575_),
    .A2(_05568_),
    .B(_05576_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11260_ (.A1(_04381_),
    .A2(_04495_),
    .A3(_04502_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11261_ (.I(_05577_),
    .Z(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11262_ (.I(_05578_),
    .Z(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11263_ (.I(_05577_),
    .Z(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11264_ (.I(_05580_),
    .Z(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11265_ (.A1(\as2650.stack[13][0] ),
    .A2(_05581_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11266_ (.A1(_05534_),
    .A2(_05579_),
    .B(_05582_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11267_ (.A1(\as2650.stack[13][1] ),
    .A2(_05581_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11268_ (.A1(_05541_),
    .A2(_05579_),
    .B(_05583_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11269_ (.A1(\as2650.stack[13][2] ),
    .A2(_05581_),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11270_ (.A1(_05543_),
    .A2(_05579_),
    .B(_05584_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11271_ (.A1(\as2650.stack[13][3] ),
    .A2(_05581_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11272_ (.A1(_05545_),
    .A2(_05579_),
    .B(_05585_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11273_ (.I(_05578_),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11274_ (.I(_05580_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11275_ (.A1(\as2650.stack[13][4] ),
    .A2(_05587_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11276_ (.A1(_05547_),
    .A2(_05586_),
    .B(_05588_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11277_ (.A1(\as2650.stack[13][5] ),
    .A2(_05587_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11278_ (.A1(_05551_),
    .A2(_05586_),
    .B(_05589_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11279_ (.A1(\as2650.stack[13][6] ),
    .A2(_05587_),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11280_ (.A1(_05553_),
    .A2(_05586_),
    .B(_05590_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11281_ (.A1(\as2650.stack[13][7] ),
    .A2(_05587_),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11282_ (.A1(_05555_),
    .A2(_05586_),
    .B(_05591_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11283_ (.I(_05578_),
    .Z(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11284_ (.I(_05580_),
    .Z(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11285_ (.A1(\as2650.stack[13][8] ),
    .A2(_05593_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11286_ (.A1(_05557_),
    .A2(_05592_),
    .B(_05594_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11287_ (.A1(\as2650.stack[13][9] ),
    .A2(_05593_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11288_ (.A1(_05561_),
    .A2(_05592_),
    .B(_05595_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11289_ (.A1(\as2650.stack[13][10] ),
    .A2(_05593_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11290_ (.A1(_05563_),
    .A2(_05592_),
    .B(_05596_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11291_ (.A1(\as2650.stack[13][11] ),
    .A2(_05593_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11292_ (.A1(_05565_),
    .A2(_05592_),
    .B(_05597_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11293_ (.I(_05578_),
    .Z(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11294_ (.I(_05580_),
    .Z(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11295_ (.A1(\as2650.stack[13][12] ),
    .A2(_05599_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11296_ (.A1(_05567_),
    .A2(_05598_),
    .B(_05600_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11297_ (.A1(\as2650.stack[13][13] ),
    .A2(_05599_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11298_ (.A1(_05571_),
    .A2(_05598_),
    .B(_05601_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11299_ (.A1(\as2650.stack[13][14] ),
    .A2(_05599_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11300_ (.A1(_05573_),
    .A2(_05598_),
    .B(_05602_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11301_ (.A1(\as2650.stack[13][15] ),
    .A2(_05599_),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11302_ (.A1(_05575_),
    .A2(_05598_),
    .B(_05603_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11303_ (.A1(_04381_),
    .A2(_04495_),
    .A3(_04657_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11304_ (.I(_05604_),
    .Z(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11305_ (.I(_05605_),
    .Z(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11306_ (.I(_05604_),
    .Z(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11307_ (.I(_05607_),
    .Z(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11308_ (.A1(\as2650.stack[12][0] ),
    .A2(_05608_),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11309_ (.A1(_05534_),
    .A2(_05606_),
    .B(_05609_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11310_ (.A1(\as2650.stack[12][1] ),
    .A2(_05608_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11311_ (.A1(_05541_),
    .A2(_05606_),
    .B(_05610_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11312_ (.A1(\as2650.stack[12][2] ),
    .A2(_05608_),
    .ZN(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11313_ (.A1(_05543_),
    .A2(_05606_),
    .B(_05611_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11314_ (.A1(\as2650.stack[12][3] ),
    .A2(_05608_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11315_ (.A1(_05545_),
    .A2(_05606_),
    .B(_05612_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11316_ (.I(_05605_),
    .Z(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11317_ (.I(_05607_),
    .Z(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11318_ (.A1(\as2650.stack[12][4] ),
    .A2(_05614_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11319_ (.A1(_05547_),
    .A2(_05613_),
    .B(_05615_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11320_ (.A1(\as2650.stack[12][5] ),
    .A2(_05614_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11321_ (.A1(_05551_),
    .A2(_05613_),
    .B(_05616_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11322_ (.A1(\as2650.stack[12][6] ),
    .A2(_05614_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11323_ (.A1(_05553_),
    .A2(_05613_),
    .B(_05617_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11324_ (.A1(\as2650.stack[12][7] ),
    .A2(_05614_),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11325_ (.A1(_05555_),
    .A2(_05613_),
    .B(_05618_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11326_ (.I(_05605_),
    .Z(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11327_ (.I(_05607_),
    .Z(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11328_ (.A1(\as2650.stack[12][8] ),
    .A2(_05620_),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11329_ (.A1(_05557_),
    .A2(_05619_),
    .B(_05621_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11330_ (.A1(\as2650.stack[12][9] ),
    .A2(_05620_),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11331_ (.A1(_05561_),
    .A2(_05619_),
    .B(_05622_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11332_ (.A1(\as2650.stack[12][10] ),
    .A2(_05620_),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11333_ (.A1(_05563_),
    .A2(_05619_),
    .B(_05623_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11334_ (.A1(\as2650.stack[12][11] ),
    .A2(_05620_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11335_ (.A1(_05565_),
    .A2(_05619_),
    .B(_05624_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11336_ (.I(_05605_),
    .Z(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11337_ (.I(_05607_),
    .Z(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11338_ (.A1(\as2650.stack[12][12] ),
    .A2(_05626_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11339_ (.A1(_05567_),
    .A2(_05625_),
    .B(_05627_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11340_ (.A1(\as2650.stack[12][13] ),
    .A2(_05626_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11341_ (.A1(_05571_),
    .A2(_05625_),
    .B(_05628_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11342_ (.A1(\as2650.stack[12][14] ),
    .A2(_05626_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11343_ (.A1(_05573_),
    .A2(_05625_),
    .B(_05629_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11344_ (.A1(\as2650.stack[12][15] ),
    .A2(_05626_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11345_ (.A1(_05575_),
    .A2(_05625_),
    .B(_05630_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11346_ (.A1(_04502_),
    .A2(_05202_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11347_ (.I(_05631_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11348_ (.I(_05632_),
    .Z(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11349_ (.I(_05631_),
    .Z(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11350_ (.I(_05634_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11351_ (.A1(\as2650.stack[9][0] ),
    .A2(_05635_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11352_ (.A1(_05534_),
    .A2(_05633_),
    .B(_05636_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11353_ (.A1(\as2650.stack[9][1] ),
    .A2(_05635_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11354_ (.A1(_05541_),
    .A2(_05633_),
    .B(_05637_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11355_ (.A1(\as2650.stack[9][2] ),
    .A2(_05635_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11356_ (.A1(_05543_),
    .A2(_05633_),
    .B(_05638_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11357_ (.A1(\as2650.stack[9][3] ),
    .A2(_05635_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11358_ (.A1(_05545_),
    .A2(_05633_),
    .B(_05639_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11359_ (.I(_05632_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11360_ (.I(_05634_),
    .Z(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11361_ (.A1(\as2650.stack[9][4] ),
    .A2(_05641_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11362_ (.A1(_05547_),
    .A2(_05640_),
    .B(_05642_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11363_ (.A1(\as2650.stack[9][5] ),
    .A2(_05641_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11364_ (.A1(_05551_),
    .A2(_05640_),
    .B(_05643_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11365_ (.A1(\as2650.stack[9][6] ),
    .A2(_05641_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11366_ (.A1(_05553_),
    .A2(_05640_),
    .B(_05644_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11367_ (.A1(\as2650.stack[9][7] ),
    .A2(_05641_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11368_ (.A1(_05555_),
    .A2(_05640_),
    .B(_05645_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11369_ (.I(_05632_),
    .Z(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11370_ (.I(_05634_),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11371_ (.A1(\as2650.stack[9][8] ),
    .A2(_05647_),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11372_ (.A1(_05557_),
    .A2(_05646_),
    .B(_05648_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11373_ (.A1(\as2650.stack[9][9] ),
    .A2(_05647_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11374_ (.A1(_05561_),
    .A2(_05646_),
    .B(_05649_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11375_ (.A1(\as2650.stack[9][10] ),
    .A2(_05647_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11376_ (.A1(_05563_),
    .A2(_05646_),
    .B(_05650_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11377_ (.A1(\as2650.stack[9][11] ),
    .A2(_05647_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11378_ (.A1(_05565_),
    .A2(_05646_),
    .B(_05651_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11379_ (.I(_05632_),
    .Z(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11380_ (.I(_05634_),
    .Z(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11381_ (.A1(\as2650.stack[9][12] ),
    .A2(_05653_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11382_ (.A1(_05567_),
    .A2(_05652_),
    .B(_05654_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11383_ (.A1(\as2650.stack[9][13] ),
    .A2(_05653_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11384_ (.A1(_05571_),
    .A2(_05652_),
    .B(_05655_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11385_ (.A1(\as2650.stack[9][14] ),
    .A2(_05653_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11386_ (.A1(_05573_),
    .A2(_05652_),
    .B(_05656_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11387_ (.A1(\as2650.stack[9][15] ),
    .A2(_05653_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11388_ (.A1(_05575_),
    .A2(_05652_),
    .B(_05657_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11389_ (.D(_00017_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11390_ (.D(_00018_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(net122));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11391_ (.D(_00019_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(net129));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11392_ (.D(_00020_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net130));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11393_ (.D(_00021_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(net131));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11394_ (.D(_00022_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11395_ (.D(_00023_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11396_ (.D(_00024_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11397_ (.D(_00025_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11398_ (.D(_00026_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11399_ (.D(_00027_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11400_ (.D(_00028_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(net123));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11401_ (.D(_00029_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(net124));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11402_ (.D(_00030_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(net125));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11403_ (.D(_00031_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(net126));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11404_ (.D(_00032_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(net127));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11405_ (.D(_00033_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(net128));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11406_ (.D(_00034_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(net106));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11407_ (.D(_00035_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(net113));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11408_ (.D(_00036_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net114));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11409_ (.D(_00037_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net115));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11410_ (.D(_00038_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net116));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11411_ (.D(_00039_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net117));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11412_ (.D(_00040_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net118));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11413_ (.D(_00041_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net119));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11414_ (.D(_00042_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(net120));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11415_ (.D(_00043_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(net121));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11416_ (.D(_00044_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(net107));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11417_ (.D(_00045_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(net108));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11418_ (.D(_00046_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net109));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11419_ (.D(_00047_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net110));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11420_ (.D(_00048_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(net111));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11421_ (.D(_00049_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(net112));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11422_ (.D(_00050_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net239));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11423_ (.D(_00051_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net159));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11424_ (.D(_00052_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net160));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11425_ (.D(_00053_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net161));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11426_ (.D(_00054_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net265));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11427_ (.D(_00055_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(net266));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11428_ (.D(_00056_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(net277));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11429_ (.D(_00057_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net288));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11430_ (.D(_00058_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net291));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11431_ (.D(_00059_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net292));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11432_ (.D(_00060_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net293));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11433_ (.D(_00061_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net294));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11434_ (.D(_00062_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net295));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11435_ (.D(_00063_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net296));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11436_ (.D(_00064_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net297));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11437_ (.D(_00065_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(net267));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11438_ (.D(_00066_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(net268));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11439_ (.D(_00067_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(net269));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11440_ (.D(_00068_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(net270));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11441_ (.D(_00069_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(net271));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11442_ (.D(_00070_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(net272));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11443_ (.D(_00071_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(net273));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11444_ (.D(_00072_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net274));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11445_ (.D(_00073_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net275));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11446_ (.D(_00074_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net276));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11447_ (.D(_00075_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net278));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11448_ (.D(_00076_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net279));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11449_ (.D(_00077_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net280));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11450_ (.D(_00078_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(net281));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11451_ (.D(_00079_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(net282));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11452_ (.D(_00080_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(net283));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11453_ (.D(_00081_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(net284));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11454_ (.D(_00082_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(net285));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11455_ (.D(_00083_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net286));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11456_ (.D(_00084_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net287));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11457_ (.D(_00085_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(net289));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11458_ (.D(_00086_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(net290));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11459_ (.D(_00087_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11460_ (.D(net366),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11461_ (.D(net363),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(wb_debug_carry));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11462_ (.D(net360),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\web_behavior[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11463_ (.D(net357),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\web_behavior[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11464_ (.D(net373),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(wb_reset_override_en));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11465_ (.D(net421),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(wb_reset_override));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11466_ (.D(_00094_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(wb_io3_test));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11467_ (.D(net396),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(net182));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11468_ (.D(_00096_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11469_ (.D(_00097_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\wb_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11470_ (.D(_00098_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\wb_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11471_ (.D(_00099_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\wb_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11472_ (.D(_00100_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\wb_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11473_ (.D(_00101_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(\wb_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11474_ (.D(_00102_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\wb_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11475_ (.D(_00103_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\wb_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11476_ (.D(_00104_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\wb_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11477_ (.D(_00105_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\wb_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11478_ (.D(_00106_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\wb_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11479_ (.D(net415),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\wb_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11480_ (.D(net418),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\wb_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11481_ (.D(net403),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\wb_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11482_ (.D(net409),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\wb_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11483_ (.D(net400),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\wb_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11484_ (.D(net385),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\wb_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11485_ (.D(net381),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\wb_counter[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11486_ (.D(net393),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\wb_counter[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11487_ (.D(net389),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\wb_counter[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11488_ (.D(net370),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\wb_counter[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11489_ (.D(net377),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\wb_counter[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11490_ (.D(_00118_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\wb_counter[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11491_ (.D(_00119_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\wb_counter[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11492_ (.D(_00120_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\wb_counter[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11493_ (.D(_00121_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\wb_counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11494_ (.D(_00122_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\wb_counter[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11495_ (.D(_00123_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\wb_counter[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11496_ (.D(_00124_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\wb_counter[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11497_ (.D(net412),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\wb_counter[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11498_ (.D(_00126_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\wb_counter[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11499_ (.D(net406),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\wb_counter[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11500_ (.D(_00128_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\wb_counter[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11501_ (.D(_00129_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(net221));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11502_ (.D(_00130_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(net228));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11503_ (.D(_00131_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(net229));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11504_ (.D(_00132_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net230));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11505_ (.D(_00133_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(net231));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11506_ (.D(_00134_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(net232));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11507_ (.D(_00135_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(net233));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11508_ (.D(_00136_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(net234));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11509_ (.D(_00137_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11510_ (.D(_00138_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.insin[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11511_ (.D(_00139_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.insin[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11512_ (.D(_00140_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.insin[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11513_ (.D(_00141_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.insin[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11514_ (.D(_00142_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.insin[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11515_ (.D(_00143_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.insin[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11516_ (.D(_00144_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.indirect_target[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11517_ (.D(_00005_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11518_ (.D(_00008_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11519_ (.D(_00009_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11520_ (.D(_00010_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.is_interrupt_cycle ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11521_ (.D(_00011_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11522_ (.D(_00012_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11523_ (.D(_00013_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11524_ (.D(_00014_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11525_ (.D(_00015_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11526_ (.D(_00016_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11527_ (.D(_00006_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11528_ (.D(_00007_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11529_ (.D(_00145_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.cpu_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11530_ (.D(_00146_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.chirp_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11531_ (.D(_00147_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.chirp_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11532_ (.D(_00148_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.chirp_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11533_ (.D(_00149_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.indirect_target[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11534_ (.D(_00150_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.indirect_target[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11535_ (.D(_00151_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.indirect_target[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11536_ (.D(_00152_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.indirect_target[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11537_ (.D(_00153_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.indirect_target[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11538_ (.D(_00154_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.indirect_target[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11539_ (.D(_00155_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.indirect_target[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11540_ (.D(_00156_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.indirect_target[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11541_ (.D(_00157_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.indirect_target[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11542_ (.D(_00158_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.indirect_target[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11543_ (.D(_00159_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.indirect_target[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11544_ (.D(_00160_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.indirect_target[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11545_ (.D(_00161_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.indirect_target[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11546_ (.D(_00162_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.indirect_target[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11547_ (.D(_00163_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.indirect_target[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11548_ (.D(_00164_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.indexed_cyc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11549_ (.D(_00165_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.indexed_cyc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11550_ (.D(_00166_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.indirect_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11551_ (.D(_00167_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.extend ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11552_ (.D(_00168_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(net213));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11553_ (.D(_00169_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11554_ (.D(_00170_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11555_ (.D(_00171_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.instruction_args_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11556_ (.D(_00172_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11557_ (.D(_00173_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.instruction_args_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11558_ (.D(_00174_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11559_ (.D(_00175_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11560_ (.D(_00176_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.instruction_args_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11561_ (.D(_00177_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11562_ (.D(_00178_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11563_ (.D(_00179_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11564_ (.D(_00180_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11565_ (.D(_00181_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11566_ (.D(_00182_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11567_ (.D(_00183_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11568_ (.D(_00184_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11569_ (.D(_00185_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\as2650.instruction_args_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11570_ (.D(_00186_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11571_ (.D(_00187_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11572_ (.D(_00188_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11573_ (.D(_00189_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11574_ (.D(_00190_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11575_ (.D(_00191_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.insin[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11576_ (.D(_00192_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11577_ (.D(_00193_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11578_ (.D(_00194_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11579_ (.D(_00195_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11580_ (.D(_00196_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11581_ (.D(_00197_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11582_ (.D(_00198_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11583_ (.D(_00199_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11584_ (.D(_00200_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11585_ (.D(_00201_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.ivectors_base[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11586_ (.D(_00202_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.ivectors_base[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11587_ (.D(_00203_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11588_ (.D(_00204_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.PC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11589_ (.D(_00205_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11590_ (.D(_00206_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11591_ (.D(_00207_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.PC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11592_ (.D(_00208_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11593_ (.D(_00209_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11594_ (.D(_00210_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11595_ (.D(_00211_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11596_ (.D(_00212_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11597_ (.D(_00213_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11598_ (.D(_00214_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11599_ (.D(_00215_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11600_ (.D(_00216_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11601_ (.D(_00217_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.debug_psl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11602_ (.D(_00218_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11603_ (.D(_00219_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11604_ (.D(_00220_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11605_ (.D(_00221_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11606_ (.D(_00222_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.debug_psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11607_ (.D(_00223_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.debug_psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11608_ (.D(_00224_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11609_ (.D(_00225_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.debug_psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11610_ (.D(_00226_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.debug_psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11611_ (.D(_00227_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.debug_psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11612_ (.D(_00228_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11613_ (.D(_00229_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11614_ (.D(_00230_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(net181));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11615_ (.D(_00231_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11616_ (.D(_00232_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.irqs_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11617_ (.D(_00233_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.irqs_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11618_ (.D(_00234_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.irqs_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11619_ (.D(_00235_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.irqs_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11620_ (.D(_00236_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.irqs_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11621_ (.D(_00237_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.irqs_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11622_ (.D(_00238_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.irqs_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11623_ (.D(_00239_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11624_ (.D(_00240_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net147));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11625_ (.D(_00241_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net148));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11626_ (.D(_00242_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net149));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11627_ (.D(_00243_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net150));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11628_ (.D(_00244_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net151));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11629_ (.D(_00245_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net152));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11630_ (.D(_00246_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net153));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11631_ (.D(_00247_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net154));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11632_ (.D(_00248_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net146));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11633_ (.D(_00249_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net140));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11634_ (.D(_00250_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net141));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11635_ (.D(_00251_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net142));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11636_ (.D(_00252_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net143));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11637_ (.D(_00253_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11638_ (.D(_00254_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(net145));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11639_ (.D(_00255_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.ext_io_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11640_ (.D(_00256_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.ext_io_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11641_ (.D(_00257_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11642_ (.D(_00258_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(net235));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11643_ (.D(_00259_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net236));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11644_ (.D(_00260_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(net222));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11645_ (.D(_00261_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(net223));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11646_ (.D(_00262_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(net224));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11647_ (.D(_00263_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net225));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11648_ (.D(_00264_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(net226));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11649_ (.D(_00265_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net227));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11650_ (.D(_00266_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11651_ (.D(_00267_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11652_ (.D(_00268_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11653_ (.D(_00269_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11654_ (.D(_00270_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11655_ (.D(_00271_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11656_ (.D(_00272_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11657_ (.D(_00273_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11658_ (.D(_00274_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11659_ (.D(_00275_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11660_ (.D(_00276_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11661_ (.D(_00277_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11662_ (.D(_00278_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11663_ (.D(_00279_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11664_ (.D(_00280_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11665_ (.D(_00281_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11666_ (.D(_00282_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11667_ (.D(_00283_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11668_ (.D(_00284_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11669_ (.D(_00285_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11670_ (.D(_00286_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11671_ (.D(_00287_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11672_ (.D(_00288_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11673_ (.D(_00289_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11674_ (.D(_00290_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11675_ (.D(_00291_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11676_ (.D(_00292_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11677_ (.D(_00293_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11678_ (.D(_00294_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11679_ (.D(_00295_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11680_ (.D(_00296_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11681_ (.D(_00297_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11682_ (.D(_00298_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11683_ (.D(_00299_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11684_ (.D(_00300_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00301_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00302_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00303_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00304_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00305_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00306_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00307_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00308_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00309_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00310_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00311_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00312_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11697_ (.D(_00313_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00314_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00315_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00316_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00317_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00318_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00319_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00320_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00321_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00322_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00323_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00324_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00325_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00326_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00327_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00328_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00329_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00330_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11715_ (.D(_00331_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00332_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00333_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00334_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00335_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00336_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00337_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00338_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00339_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11724_ (.D(_00340_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00341_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00342_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00343_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00344_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00345_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00346_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00347_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00348_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00349_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00350_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00351_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00352_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00353_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00354_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00355_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00356_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00357_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00358_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00359_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00360_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00361_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00362_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00363_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00364_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00365_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00366_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00367_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00368_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00369_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00370_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00371_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00372_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00373_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00374_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00375_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00376_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11761_ (.D(_00377_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11762_ (.D(_00378_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11763_ (.D(_00379_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11764_ (.D(_00380_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11765_ (.D(_00381_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00382_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11767_ (.D(_00383_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11768_ (.D(_00384_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00385_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00386_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00387_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00388_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00389_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00390_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00391_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00392_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00393_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00394_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00395_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00396_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00397_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00398_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00399_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00400_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00401_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00402_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00403_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00404_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00405_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00406_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00407_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00408_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00409_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00410_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00411_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00412_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00413_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00414_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00415_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00416_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00417_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00418_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00419_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00420_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00421_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00422_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00423_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00424_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00425_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00426_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00427_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11812_ (.D(_00428_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11813_ (.D(_00429_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11814_ (.D(_00430_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00431_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11816_ (.D(_00432_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11817_ (.D(_00433_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11818_ (.D(_00434_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00435_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11820_ (.D(_00436_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11821_ (.D(_00437_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00438_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00439_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00440_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00441_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00442_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.chirpchar[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00443_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00444_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00445_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11830_ (.D(_00446_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00447_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00448_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00449_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00450_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00451_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00452_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00453_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00454_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00455_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11840_ (.D(_00456_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11841_ (.D(_00457_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11842_ (.D(_00458_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00459_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00460_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00461_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00462_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00463_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11848_ (.D(_00464_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11849_ (.D(_00465_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00466_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00467_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00468_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00469_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00470_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00471_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00472_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00473_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00474_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11859_ (.D(_00475_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00476_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00477_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11862_ (.D(_00478_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00479_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00480_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00481_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00482_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00483_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00484_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00485_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00486_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00487_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00488_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11873_ (.D(_00489_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11874_ (.D(_00490_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11875_ (.D(_00491_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11876_ (.D(_00492_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11877_ (.D(_00493_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00494_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00495_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00496_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00497_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00498_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00499_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00500_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00501_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00502_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00503_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00504_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11889_ (.D(_00505_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11890_ (.D(_00506_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11891_ (.D(_00507_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11892_ (.D(_00508_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11893_ (.D(_00509_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.regs[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11894_ (.D(_00510_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11895_ (.D(_00511_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11896_ (.D(_00512_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11897_ (.D(_00513_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11898_ (.D(_00514_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11899_ (.D(_00000_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.chirpchar[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00001_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.chirpchar[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11901_ (.D(_00002_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.chirpchar[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00003_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.chirpchar[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00004_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.chirpchar[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00515_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.chirpchar[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00516_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11906_ (.D(_00517_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11907_ (.D(_00518_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11908_ (.D(_00519_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11909_ (.D(_00520_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00521_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00522_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11912_ (.D(_00523_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00524_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00525_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11915_ (.D(_00526_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11916_ (.D(_00527_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11917_ (.D(_00528_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11918_ (.D(_00529_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11919_ (.D(_00530_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00531_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00532_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00533_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00534_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11924_ (.D(_00535_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11925_ (.D(_00536_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11926_ (.D(_00537_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11927_ (.D(_00538_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11928_ (.D(_00539_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11929_ (.D(_00540_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11930_ (.D(_00541_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00542_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00543_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00544_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00545_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00546_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11936_ (.D(_00547_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11937_ (.D(_00548_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00549_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11939_ (.D(_00550_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11940_ (.D(_00551_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11941_ (.D(_00552_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11942_ (.D(_00553_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_00554_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11944_ (.D(_00555_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11945_ (.D(_00556_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_00557_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_00558_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11948_ (.D(_00559_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11949_ (.D(_00560_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11950_ (.D(_00561_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11951_ (.D(_00562_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_00563_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_00564_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11954_ (.D(_00565_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_00566_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11956_ (.D(_00567_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11957_ (.D(_00568_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_00569_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_00570_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11960_ (.D(_00571_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11961_ (.D(_00572_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11962_ (.D(_00573_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11963_ (.D(_00574_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11964_ (.D(_00575_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_00576_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_00577_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_00578_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_00579_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11969_ (.D(_00580_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_00581_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11971_ (.D(_00582_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11972_ (.D(_00583_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11973_ (.D(_00584_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11974_ (.D(_00585_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11975_ (.D(_00586_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11976_ (.D(_00587_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12015_ (.I(net306),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12016_ (.I(net306),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12017_ (.I(net306),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12018_ (.I(net307),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12019_ (.I(net307),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12020_ (.I(net307),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12021_ (.I(net308),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12022_ (.I(net306),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12023_ (.I(net305),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12024_ (.I(net304),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12025_ (.I(net303),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12026_ (.I(net302),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12027_ (.I(net301),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12028_ (.I(net300),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12029_ (.I(net299),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12030_ (.I(net298),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_110_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_118_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_128_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_129_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_130_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_132_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_135_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_137_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_138_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_139_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_142_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_144_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_145_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_84_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_90_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout306 (.I(net307),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout307 (.I(net164),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout308 (.I(net164),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(net453),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold100 (.I(wbs_dat_i[15]),
    .Z(net449));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold101 (.I(wbs_dat_i[17]),
    .Z(net450));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold102 (.I(wbs_dat_i[1]),
    .Z(net451));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold103 (.I(wbs_dat_i[13]),
    .Z(net452));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold104 (.I(wbs_dat_i[2]),
    .Z(net453));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold105 (.I(wbs_dat_i[22]),
    .Z(net454));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold106 (.I(wbs_dat_i[11]),
    .Z(net455));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold107 (.I(wbs_dat_i[0]),
    .Z(net456));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold108 (.I(wbs_dat_i[12]),
    .Z(net457));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold109 (.I(wbs_dat_i[3]),
    .Z(net458));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(_01988_),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold110 (.I(wbs_dat_i[21]),
    .Z(net459));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold111 (.I(wbs_dat_i[6]),
    .Z(net460));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold112 (.I(wbs_dat_i[25]),
    .Z(net461));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold113 (.I(wbs_dat_i[23]),
    .Z(net462));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold114 (.I(wbs_dat_i[9]),
    .Z(net463));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold115 (.I(wbs_dat_i[10]),
    .Z(net464));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold116 (.I(wbs_dat_i[26]),
    .Z(net465));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold117 (.I(wbs_dat_i[4]),
    .Z(net466));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold118 (.I(wbs_dat_i[24]),
    .Z(net467));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold119 (.I(wbs_dat_i[18]),
    .Z(net468));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(_00090_),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold120 (.I(wbs_dat_i[30]),
    .Z(net469));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold121 (.I(wbs_dat_i[20]),
    .Z(net470));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold122 (.I(wbs_dat_i[27]),
    .Z(net471));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold123 (.I(wbs_dat_i[5]),
    .Z(net472));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold124 (.I(wbs_adr_i[22]),
    .Z(net473));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold125 (.I(wbs_dat_i[19]),
    .Z(net474));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold126 (.I(wbs_adr_i[19]),
    .Z(net475));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold127 (.I(_01764_),
    .Z(net476));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold128 (.I(wbs_dat_i[28]),
    .Z(net477));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold129 (.I(wbs_adr_i[20]),
    .Z(net478));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(net451),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold130 (.I(wbs_dat_i[16]),
    .Z(net479));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(_01984_),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(_00089_),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(net456),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(_01982_),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(_00088_),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(net474),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(net82),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(_02081_),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(_00116_),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(net466),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(_01992_),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(_00092_),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(net470),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(net84),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(_02086_),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(_00117_),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(net479),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(net79),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(_02070_),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(_00113_),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(net449),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(net78),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(_02066_),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(_00112_),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(net468),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(net81),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(_02078_),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(_00115_),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(net450),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(net80),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(_02075_),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(_00114_),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(net448),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(_01997_),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(_00095_),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(net446),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(net77),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(_02061_),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(_00111_),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(net457),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(_02054_),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(_00109_),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(net469),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(_02125_),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(_00127_),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(net452),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(_02058_),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(_00110_),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(net477),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(_02118_),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(_00125_),
    .Z(net412));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(net464),
    .Z(net413));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(_02045_),
    .Z(net414));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(_00107_),
    .Z(net415));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(net455),
    .Z(net416));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(_02048_),
    .Z(net417));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(net458),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(_00108_),
    .Z(net418));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(net472),
    .Z(net419));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(_01994_),
    .Z(net420));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(_00093_),
    .Z(net421));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(net473),
    .Z(net422));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(net443),
    .Z(net423));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(net444),
    .Z(net424));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(net445),
    .Z(net425));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(net447),
    .Z(net426));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold79 (.I(net69),
    .Z(net427));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(_01990_),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(net478),
    .Z(net428));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(net454),
    .Z(net429));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(net459),
    .Z(net430));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(net461),
    .Z(net431));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(net462),
    .Z(net432));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(net460),
    .Z(net433));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(net463),
    .Z(net434));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(net467),
    .Z(net435));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(net475),
    .Z(net436));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold89 (.I(_01729_),
    .Z(net437));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(_00091_),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(net465),
    .Z(net438));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(net471),
    .Z(net439));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(wbs_cyc_i),
    .Z(net440));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(_01664_),
    .Z(net441));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold94 (.I(wbs_dat_i[29]),
    .Z(net443));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold95 (.I(wbs_dat_i[31]),
    .Z(net444));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold96 (.I(wbs_dat_i[8]),
    .Z(net445));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold97 (.I(wbs_dat_i[14]),
    .Z(net446));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold98 (.I(wbs_adr_i[21]),
    .Z(net447));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold99 (.I(wbs_dat_i[7]),
    .Z(net448));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(bus_in_gpios[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(bus_in_serial_ports[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input100 (.I(net433),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input101 (.I(net394),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input102 (.I(net425),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input103 (.I(net434),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input104 (.I(wbs_stb_i),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input105 (.I(wbs_we_i),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(bus_in_serial_ports[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input12 (.I(bus_in_serial_ports[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(bus_in_serial_ports[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(bus_in_serial_ports[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(bus_in_serial_ports[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(bus_in_serial_ports[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(bus_in_sid[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(bus_in_sid[1]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(bus_in_sid[2]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(bus_in_gpios[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(bus_in_sid[3]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(bus_in_sid[4]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(bus_in_sid[5]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(bus_in_sid[6]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(bus_in_sid[7]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(bus_in_timers[0]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(bus_in_timers[1]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(bus_in_timers[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(bus_in_timers[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(bus_in_timers[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(bus_in_gpios[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(bus_in_timers[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(bus_in_timers[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(bus_in_timers[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input33 (.I(io_in[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input34 (.I(io_in[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input35 (.I(io_in[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(io_in[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input37 (.I(io_in[4]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(io_in[5]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(io_in[6]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(bus_in_gpios[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(io_in[7]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(io_in[8]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input42 (.I(io_in[9]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(irqs[0]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input44 (.I(irqs[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input45 (.I(irqs[2]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input46 (.I(irqs[3]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(irqs[4]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input48 (.I(irqs[5]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(irqs[6]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(bus_in_gpios[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input50 (.I(ram_bus_in[0]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(ram_bus_in[1]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(ram_bus_in[2]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(ram_bus_in[3]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(ram_bus_in[4]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(ram_bus_in[5]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(ram_bus_in[6]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(ram_bus_in[7]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input58 (.I(rom_bus_in[0]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input59 (.I(rom_bus_in[1]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(bus_in_gpios[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input60 (.I(rom_bus_in[2]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input61 (.I(rom_bus_in[3]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input62 (.I(rom_bus_in[4]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input63 (.I(rom_bus_in[5]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input64 (.I(rom_bus_in[6]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input65 (.I(rom_bus_in[7]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input66 (.I(wb_rst_i),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input67 (.I(net436),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input68 (.I(net428),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input69 (.I(net426),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(bus_in_gpios[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input70 (.I(net422),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(net440),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input72 (.I(net364),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input73 (.I(net413),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input74 (.I(net416),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input75 (.I(net401),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(net407),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(net397),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(net382),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(net378),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(bus_in_gpios[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(net390),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(net386),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input82 (.I(net367),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input83 (.I(net361),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input84 (.I(net374),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input85 (.I(net430),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(net429),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(net432),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(net435),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input89 (.I(net431),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(bus_in_serial_ports[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input90 (.I(net438),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input91 (.I(net439),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input92 (.I(net410),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input93 (.I(net423),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input94 (.I(net358),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input95 (.I(net404),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input96 (.I(net424),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input97 (.I(net355),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input98 (.I(net371),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input99 (.I(net419),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap309 (.I(_01492_),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(RAM_end_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(RAM_end_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(RAM_end_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(RAM_end_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(RAM_end_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(RAM_end_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(RAM_end_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(RAM_end_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(RAM_end_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(RAM_end_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(RAM_end_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(RAM_end_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(RAM_end_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(RAM_end_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(RAM_end_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(RAM_end_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(RAM_start_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(RAM_start_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output124 (.I(net124),
    .Z(RAM_start_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output125 (.I(net125),
    .Z(RAM_start_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output126 (.I(net126),
    .Z(RAM_start_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output127 (.I(net127),
    .Z(RAM_start_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output128 (.I(net128),
    .Z(RAM_start_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output129 (.I(net129),
    .Z(RAM_start_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output130 (.I(net130),
    .Z(RAM_start_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output131 (.I(net131),
    .Z(RAM_start_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output132 (.I(net132),
    .Z(RAM_start_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output133 (.I(net133),
    .Z(RAM_start_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output134 (.I(net134),
    .Z(RAM_start_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output135 (.I(net135),
    .Z(RAM_start_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output136 (.I(net136),
    .Z(RAM_start_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output137 (.I(net137),
    .Z(RAM_start_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output138 (.I(net138),
    .Z(WEb_raw));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output139 (.I(net139),
    .Z(boot_rom_en));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output140 (.I(net140),
    .Z(bus_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output141 (.I(net141),
    .Z(bus_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output142 (.I(net142),
    .Z(bus_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output143 (.I(net143),
    .Z(bus_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output144 (.I(net144),
    .Z(bus_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output145 (.I(net145),
    .Z(bus_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output146 (.I(net146),
    .Z(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output147 (.I(net147),
    .Z(bus_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output148 (.I(net148),
    .Z(bus_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output149 (.I(net149),
    .Z(bus_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output150 (.I(net150),
    .Z(bus_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output151 (.I(net151),
    .Z(bus_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output152 (.I(net152),
    .Z(bus_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output153 (.I(net153),
    .Z(bus_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output154 (.I(net154),
    .Z(bus_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output155 (.I(net155),
    .Z(bus_we_gpios));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output156 (.I(net156),
    .Z(bus_we_serial_ports));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output157 (.I(net157),
    .Z(bus_we_sid));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output158 (.I(net158),
    .Z(bus_we_timers));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output159 (.I(net159),
    .Z(cs_port[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output160 (.I(net160),
    .Z(cs_port[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output161 (.I(net161),
    .Z(cs_port[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output162 (.I(net162),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output163 (.I(net163),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output164 (.I(net308),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output165 (.I(net165),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output166 (.I(net166),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output167 (.I(net167),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output168 (.I(net168),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output169 (.I(net169),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output170 (.I(net170),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output171 (.I(net300),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output172 (.I(net299),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output173 (.I(net298),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output174 (.I(net174),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output175 (.I(net175),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output176 (.I(net176),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output177 (.I(net177),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output178 (.I(net178),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output179 (.I(net179),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output180 (.I(net180),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output181 (.I(net181),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output182 (.I(net182),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output183 (.I(net305),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output184 (.I(net304),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output185 (.I(net303),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output186 (.I(net302),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output187 (.I(net301),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output188 (.I(net188),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output189 (.I(net189),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output190 (.I(net190),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output191 (.I(net191),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output192 (.I(net192),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output193 (.I(net193),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output194 (.I(net194),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output195 (.I(net195),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output196 (.I(net196),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output197 (.I(net197),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output198 (.I(net198),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output199 (.I(net199),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output200 (.I(net200),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output201 (.I(net201),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output202 (.I(net202),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output203 (.I(net203),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output204 (.I(net204),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output205 (.I(net205),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output206 (.I(net206),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output207 (.I(net207),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output208 (.I(net208),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output209 (.I(net209),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output210 (.I(net210),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output211 (.I(net211),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output212 (.I(net212),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output213 (.I(net213),
    .Z(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output214 (.I(net214),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output215 (.I(net215),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output216 (.I(net216),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output217 (.I(net217),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output218 (.I(net218),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output219 (.I(net219),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output220 (.I(net220),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output221 (.I(net221),
    .Z(last_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output222 (.I(net222),
    .Z(last_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output223 (.I(net223),
    .Z(last_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output224 (.I(net224),
    .Z(last_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output225 (.I(net225),
    .Z(last_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output226 (.I(net226),
    .Z(last_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output227 (.I(net227),
    .Z(last_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output228 (.I(net228),
    .Z(last_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output229 (.I(net229),
    .Z(last_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output230 (.I(net230),
    .Z(last_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output231 (.I(net231),
    .Z(last_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output232 (.I(net232),
    .Z(last_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output233 (.I(net233),
    .Z(last_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output234 (.I(net234),
    .Z(last_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output235 (.I(net235),
    .Z(last_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output236 (.I(net236),
    .Z(last_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output237 (.I(net237),
    .Z(le_hi_act));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output238 (.I(net238),
    .Z(le_lo_act));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output239 (.I(net239),
    .Z(ram_enabled));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output240 (.I(net240),
    .Z(requested_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output241 (.I(net241),
    .Z(requested_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output242 (.I(net242),
    .Z(requested_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output243 (.I(net243),
    .Z(requested_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output244 (.I(net244),
    .Z(requested_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output245 (.I(net245),
    .Z(requested_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output246 (.I(net246),
    .Z(requested_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output247 (.I(net247),
    .Z(requested_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output248 (.I(net248),
    .Z(requested_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output249 (.I(net249),
    .Z(requested_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output250 (.I(net250),
    .Z(requested_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output251 (.I(net251),
    .Z(requested_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output252 (.I(net252),
    .Z(requested_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output253 (.I(net253),
    .Z(requested_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output254 (.I(net254),
    .Z(requested_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output255 (.I(net255),
    .Z(requested_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output256 (.I(net350),
    .Z(reset_out));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output257 (.I(net257),
    .Z(rom_bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output258 (.I(net258),
    .Z(rom_bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output259 (.I(net259),
    .Z(rom_bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output260 (.I(net260),
    .Z(rom_bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output261 (.I(net261),
    .Z(rom_bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output262 (.I(net262),
    .Z(rom_bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output263 (.I(net263),
    .Z(rom_bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output264 (.I(net264),
    .Z(rom_bus_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output265 (.I(net265),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output266 (.I(net266),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output267 (.I(net267),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output268 (.I(net268),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output269 (.I(net269),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output270 (.I(net270),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output271 (.I(net271),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output272 (.I(net272),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output273 (.I(net273),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output274 (.I(net274),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output275 (.I(net275),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output276 (.I(net276),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output277 (.I(net277),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output278 (.I(net278),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output279 (.I(net279),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output280 (.I(net280),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output281 (.I(net281),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output282 (.I(net282),
    .Z(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output283 (.I(net283),
    .Z(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output284 (.I(net284),
    .Z(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output285 (.I(net285),
    .Z(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output286 (.I(net286),
    .Z(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output287 (.I(net287),
    .Z(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output288 (.I(net288),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output289 (.I(net289),
    .Z(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output290 (.I(net290),
    .Z(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output291 (.I(net291),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output292 (.I(net292),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output293 (.I(net293),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output294 (.I(net294),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output295 (.I(net295),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output296 (.I(net296),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output297 (.I(net297),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer1 (.I(net354),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 rebuffer2 (.I(net256),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer3 (.I(_04038_),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer4 (.I(_04038_),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer5 (.I(_00681_),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer6 (.I(net442),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 rebuffer7 (.I(_00842_),
    .Z(net442));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire298 (.I(net173),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire299 (.I(net172),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire300 (.I(net171),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire301 (.I(net187),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire302 (.I(net186),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire303 (.I(net185),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire304 (.I(net184),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire305 (.I(net183),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_310 (.ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_311 (.ZN(net311));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_312 (.ZN(net312));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_313 (.ZN(net313));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_314 (.ZN(net314));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_315 (.ZN(net315));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_316 (.ZN(net316));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_317 (.ZN(net317));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_318 (.ZN(net318));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_319 (.ZN(net319));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_320 (.ZN(net320));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_321 (.ZN(net321));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_322 (.ZN(net322));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_323 (.ZN(net323));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_324 (.ZN(net324));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_325 (.ZN(net325));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_326 (.ZN(net326));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_327 (.ZN(net327));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_328 (.ZN(net328));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_329 (.ZN(net329));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_330 (.ZN(net330));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_331 (.Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_332 (.Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_333 (.Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_334 (.Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_335 (.Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_336 (.Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_337 (.Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_338 (.Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_339 (.Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_340 (.Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_341 (.Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_342 (.Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_343 (.Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_344 (.Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_345 (.Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_346 (.Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_347 (.Z(net347));
 assign io_oeb[0] = net331;
 assign io_oeb[13] = net312;
 assign io_oeb[14] = net313;
 assign io_oeb[15] = net314;
 assign io_oeb[16] = net315;
 assign io_oeb[17] = net316;
 assign io_oeb[18] = net317;
 assign io_oeb[1] = net310;
 assign io_oeb[2] = net311;
 assign io_oeb[4] = net332;
 assign io_out[0] = net318;
 assign io_out[4] = net319;
 assign irq[0] = net320;
 assign irq[1] = net321;
 assign irq[2] = net322;
 assign la_data_out[33] = net333;
 assign la_data_out[34] = net334;
 assign la_data_out[35] = net335;
 assign la_data_out[36] = net336;
 assign la_data_out[37] = net337;
 assign la_data_out[38] = net338;
 assign la_data_out[39] = net339;
 assign la_data_out[40] = net340;
 assign la_data_out[41] = net323;
 assign la_data_out[42] = net324;
 assign la_data_out[43] = net325;
 assign la_data_out[44] = net326;
 assign la_data_out[45] = net327;
 assign la_data_out[46] = net328;
 assign la_data_out[47] = net329;
 assign la_data_out[48] = net330;
 assign la_data_out[49] = net341;
 assign la_data_out[50] = net342;
 assign la_data_out[51] = net343;
 assign la_data_out[52] = net344;
 assign la_data_out[53] = net345;
 assign la_data_out[54] = net346;
 assign la_data_out[55] = net347;
endmodule

