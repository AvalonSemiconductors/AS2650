// This is the unpowered netlist.
module wrapped_as2650 (WEb_ram,
    boot_rom_en,
    bus_cyc,
    bus_we_gpios,
    bus_we_serial_ports,
    bus_we_sid,
    bus_we_timers,
    le_hi_act,
    le_lo_act,
    ram_enabled,
    reset_out,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    RAM_end_addr,
    RAM_start_addr,
    bus_addr,
    bus_data_out,
    bus_in_gpios,
    bus_in_serial_ports,
    bus_in_sid,
    bus_in_timers,
    cs_port,
    io_in,
    io_oeb,
    io_out,
    irq,
    irqs,
    la_data_out,
    last_addr,
    ram_bus_in,
    requested_addr,
    rom_bus_in,
    rom_bus_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output WEb_ram;
 output boot_rom_en;
 output bus_cyc;
 output bus_we_gpios;
 output bus_we_serial_ports;
 output bus_we_sid;
 output bus_we_timers;
 output le_hi_act;
 output le_lo_act;
 output ram_enabled;
 output reset_out;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [15:0] RAM_end_addr;
 output [15:0] RAM_start_addr;
 output [5:0] bus_addr;
 output [7:0] bus_data_out;
 input [7:0] bus_in_gpios;
 input [7:0] bus_in_serial_ports;
 input [7:0] bus_in_sid;
 input [7:0] bus_in_timers;
 output [2:0] cs_port;
 input [18:0] io_in;
 output [18:0] io_oeb;
 output [18:0] io_out;
 output [2:0] irq;
 input [6:0] irqs;
 output [55:0] la_data_out;
 output [15:0] last_addr;
 input [7:0] ram_bus_in;
 output [15:0] requested_addr;
 input [7:0] rom_bus_in;
 output [7:0] rom_bus_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire net328;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net307;
 wire net308;
 wire net329;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire \as2650.PC[0] ;
 wire \as2650.PC[10] ;
 wire \as2650.PC[11] ;
 wire \as2650.PC[12] ;
 wire \as2650.PC[1] ;
 wire \as2650.PC[2] ;
 wire \as2650.PC[3] ;
 wire \as2650.PC[4] ;
 wire \as2650.PC[5] ;
 wire \as2650.PC[6] ;
 wire \as2650.PC[7] ;
 wire \as2650.PC[8] ;
 wire \as2650.PC[9] ;
 wire \as2650.chirp_ptr[0] ;
 wire \as2650.chirp_ptr[1] ;
 wire \as2650.chirp_ptr[2] ;
 wire \as2650.chirpchar[0] ;
 wire \as2650.chirpchar[1] ;
 wire \as2650.chirpchar[2] ;
 wire \as2650.chirpchar[3] ;
 wire \as2650.chirpchar[4] ;
 wire \as2650.chirpchar[5] ;
 wire \as2650.chirpchar[6] ;
 wire \as2650.cpu_hidden_rom_enable ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[10] ;
 wire \as2650.cycle[11] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.cycle[8] ;
 wire \as2650.cycle[9] ;
 wire \as2650.debug_psl[0] ;
 wire \as2650.debug_psl[1] ;
 wire \as2650.debug_psl[2] ;
 wire \as2650.debug_psl[3] ;
 wire \as2650.debug_psl[4] ;
 wire \as2650.debug_psl[5] ;
 wire \as2650.debug_psl[6] ;
 wire \as2650.debug_psl[7] ;
 wire \as2650.debug_psu[0] ;
 wire \as2650.debug_psu[1] ;
 wire \as2650.debug_psu[2] ;
 wire \as2650.debug_psu[3] ;
 wire \as2650.debug_psu[4] ;
 wire \as2650.debug_psu[5] ;
 wire \as2650.debug_psu[7] ;
 wire \as2650.ext_io_addr[6] ;
 wire \as2650.ext_io_addr[7] ;
 wire \as2650.extend ;
 wire \as2650.indexed_cyc[0] ;
 wire \as2650.indexed_cyc[1] ;
 wire \as2650.indirect_cyc ;
 wire \as2650.indirect_target[0] ;
 wire \as2650.indirect_target[10] ;
 wire \as2650.indirect_target[11] ;
 wire \as2650.indirect_target[12] ;
 wire \as2650.indirect_target[13] ;
 wire \as2650.indirect_target[14] ;
 wire \as2650.indirect_target[15] ;
 wire \as2650.indirect_target[1] ;
 wire \as2650.indirect_target[2] ;
 wire \as2650.indirect_target[3] ;
 wire \as2650.indirect_target[4] ;
 wire \as2650.indirect_target[5] ;
 wire \as2650.indirect_target[6] ;
 wire \as2650.indirect_target[7] ;
 wire \as2650.indirect_target[8] ;
 wire \as2650.indirect_target[9] ;
 wire \as2650.insin[0] ;
 wire \as2650.insin[1] ;
 wire \as2650.insin[2] ;
 wire \as2650.insin[3] ;
 wire \as2650.insin[4] ;
 wire \as2650.insin[5] ;
 wire \as2650.insin[6] ;
 wire \as2650.insin[7] ;
 wire \as2650.instruction_args_latch[0] ;
 wire \as2650.instruction_args_latch[10] ;
 wire \as2650.instruction_args_latch[11] ;
 wire \as2650.instruction_args_latch[12] ;
 wire \as2650.instruction_args_latch[13] ;
 wire \as2650.instruction_args_latch[14] ;
 wire \as2650.instruction_args_latch[15] ;
 wire \as2650.instruction_args_latch[1] ;
 wire \as2650.instruction_args_latch[2] ;
 wire \as2650.instruction_args_latch[3] ;
 wire \as2650.instruction_args_latch[4] ;
 wire \as2650.instruction_args_latch[5] ;
 wire \as2650.instruction_args_latch[6] ;
 wire \as2650.instruction_args_latch[7] ;
 wire \as2650.instruction_args_latch[8] ;
 wire \as2650.instruction_args_latch[9] ;
 wire \as2650.io_bus_we ;
 wire \as2650.irqs_latch[1] ;
 wire \as2650.irqs_latch[2] ;
 wire \as2650.irqs_latch[3] ;
 wire \as2650.irqs_latch[4] ;
 wire \as2650.irqs_latch[5] ;
 wire \as2650.irqs_latch[6] ;
 wire \as2650.irqs_latch[7] ;
 wire \as2650.is_interrupt_cycle ;
 wire \as2650.ivectors_base[0] ;
 wire \as2650.ivectors_base[10] ;
 wire \as2650.ivectors_base[11] ;
 wire \as2650.ivectors_base[1] ;
 wire \as2650.ivectors_base[2] ;
 wire \as2650.ivectors_base[3] ;
 wire \as2650.ivectors_base[4] ;
 wire \as2650.ivectors_base[5] ;
 wire \as2650.ivectors_base[6] ;
 wire \as2650.ivectors_base[7] ;
 wire \as2650.ivectors_base[8] ;
 wire \as2650.ivectors_base[9] ;
 wire \as2650.page_reg[0] ;
 wire \as2650.page_reg[1] ;
 wire \as2650.page_reg[2] ;
 wire \as2650.regs[0][0] ;
 wire \as2650.regs[0][1] ;
 wire \as2650.regs[0][2] ;
 wire \as2650.regs[0][3] ;
 wire \as2650.regs[0][4] ;
 wire \as2650.regs[0][5] ;
 wire \as2650.regs[0][6] ;
 wire \as2650.regs[0][7] ;
 wire \as2650.regs[1][0] ;
 wire \as2650.regs[1][1] ;
 wire \as2650.regs[1][2] ;
 wire \as2650.regs[1][3] ;
 wire \as2650.regs[1][4] ;
 wire \as2650.regs[1][5] ;
 wire \as2650.regs[1][6] ;
 wire \as2650.regs[1][7] ;
 wire \as2650.regs[2][0] ;
 wire \as2650.regs[2][1] ;
 wire \as2650.regs[2][2] ;
 wire \as2650.regs[2][3] ;
 wire \as2650.regs[2][4] ;
 wire \as2650.regs[2][5] ;
 wire \as2650.regs[2][6] ;
 wire \as2650.regs[2][7] ;
 wire \as2650.regs[3][0] ;
 wire \as2650.regs[3][1] ;
 wire \as2650.regs[3][2] ;
 wire \as2650.regs[3][3] ;
 wire \as2650.regs[3][4] ;
 wire \as2650.regs[3][5] ;
 wire \as2650.regs[3][6] ;
 wire \as2650.regs[3][7] ;
 wire \as2650.regs[4][0] ;
 wire \as2650.regs[4][1] ;
 wire \as2650.regs[4][2] ;
 wire \as2650.regs[4][3] ;
 wire \as2650.regs[4][4] ;
 wire \as2650.regs[4][5] ;
 wire \as2650.regs[4][6] ;
 wire \as2650.regs[4][7] ;
 wire \as2650.regs[5][0] ;
 wire \as2650.regs[5][1] ;
 wire \as2650.regs[5][2] ;
 wire \as2650.regs[5][3] ;
 wire \as2650.regs[5][4] ;
 wire \as2650.regs[5][5] ;
 wire \as2650.regs[5][6] ;
 wire \as2650.regs[5][7] ;
 wire \as2650.regs[6][0] ;
 wire \as2650.regs[6][1] ;
 wire \as2650.regs[6][2] ;
 wire \as2650.regs[6][3] ;
 wire \as2650.regs[6][4] ;
 wire \as2650.regs[6][5] ;
 wire \as2650.regs[6][6] ;
 wire \as2650.regs[6][7] ;
 wire \as2650.regs[7][0] ;
 wire \as2650.regs[7][1] ;
 wire \as2650.regs[7][2] ;
 wire \as2650.regs[7][3] ;
 wire \as2650.regs[7][4] ;
 wire \as2650.regs[7][5] ;
 wire \as2650.regs[7][6] ;
 wire \as2650.regs[7][7] ;
 wire \as2650.relative_cyc ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][15] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[10][0] ;
 wire \as2650.stack[10][10] ;
 wire \as2650.stack[10][11] ;
 wire \as2650.stack[10][12] ;
 wire \as2650.stack[10][13] ;
 wire \as2650.stack[10][14] ;
 wire \as2650.stack[10][15] ;
 wire \as2650.stack[10][1] ;
 wire \as2650.stack[10][2] ;
 wire \as2650.stack[10][3] ;
 wire \as2650.stack[10][4] ;
 wire \as2650.stack[10][5] ;
 wire \as2650.stack[10][6] ;
 wire \as2650.stack[10][7] ;
 wire \as2650.stack[10][8] ;
 wire \as2650.stack[10][9] ;
 wire \as2650.stack[11][0] ;
 wire \as2650.stack[11][10] ;
 wire \as2650.stack[11][11] ;
 wire \as2650.stack[11][12] ;
 wire \as2650.stack[11][13] ;
 wire \as2650.stack[11][14] ;
 wire \as2650.stack[11][15] ;
 wire \as2650.stack[11][1] ;
 wire \as2650.stack[11][2] ;
 wire \as2650.stack[11][3] ;
 wire \as2650.stack[11][4] ;
 wire \as2650.stack[11][5] ;
 wire \as2650.stack[11][6] ;
 wire \as2650.stack[11][7] ;
 wire \as2650.stack[11][8] ;
 wire \as2650.stack[11][9] ;
 wire \as2650.stack[12][0] ;
 wire \as2650.stack[12][10] ;
 wire \as2650.stack[12][11] ;
 wire \as2650.stack[12][12] ;
 wire \as2650.stack[12][13] ;
 wire \as2650.stack[12][14] ;
 wire \as2650.stack[12][15] ;
 wire \as2650.stack[12][1] ;
 wire \as2650.stack[12][2] ;
 wire \as2650.stack[12][3] ;
 wire \as2650.stack[12][4] ;
 wire \as2650.stack[12][5] ;
 wire \as2650.stack[12][6] ;
 wire \as2650.stack[12][7] ;
 wire \as2650.stack[12][8] ;
 wire \as2650.stack[12][9] ;
 wire \as2650.stack[13][0] ;
 wire \as2650.stack[13][10] ;
 wire \as2650.stack[13][11] ;
 wire \as2650.stack[13][12] ;
 wire \as2650.stack[13][13] ;
 wire \as2650.stack[13][14] ;
 wire \as2650.stack[13][15] ;
 wire \as2650.stack[13][1] ;
 wire \as2650.stack[13][2] ;
 wire \as2650.stack[13][3] ;
 wire \as2650.stack[13][4] ;
 wire \as2650.stack[13][5] ;
 wire \as2650.stack[13][6] ;
 wire \as2650.stack[13][7] ;
 wire \as2650.stack[13][8] ;
 wire \as2650.stack[13][9] ;
 wire \as2650.stack[14][0] ;
 wire \as2650.stack[14][10] ;
 wire \as2650.stack[14][11] ;
 wire \as2650.stack[14][12] ;
 wire \as2650.stack[14][13] ;
 wire \as2650.stack[14][14] ;
 wire \as2650.stack[14][15] ;
 wire \as2650.stack[14][1] ;
 wire \as2650.stack[14][2] ;
 wire \as2650.stack[14][3] ;
 wire \as2650.stack[14][4] ;
 wire \as2650.stack[14][5] ;
 wire \as2650.stack[14][6] ;
 wire \as2650.stack[14][7] ;
 wire \as2650.stack[14][8] ;
 wire \as2650.stack[14][9] ;
 wire \as2650.stack[15][0] ;
 wire \as2650.stack[15][10] ;
 wire \as2650.stack[15][11] ;
 wire \as2650.stack[15][12] ;
 wire \as2650.stack[15][13] ;
 wire \as2650.stack[15][14] ;
 wire \as2650.stack[15][15] ;
 wire \as2650.stack[15][1] ;
 wire \as2650.stack[15][2] ;
 wire \as2650.stack[15][3] ;
 wire \as2650.stack[15][4] ;
 wire \as2650.stack[15][5] ;
 wire \as2650.stack[15][6] ;
 wire \as2650.stack[15][7] ;
 wire \as2650.stack[15][8] ;
 wire \as2650.stack[15][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][15] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][15] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][15] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][15] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][15] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][15] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][15] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack[8][0] ;
 wire \as2650.stack[8][10] ;
 wire \as2650.stack[8][11] ;
 wire \as2650.stack[8][12] ;
 wire \as2650.stack[8][13] ;
 wire \as2650.stack[8][14] ;
 wire \as2650.stack[8][15] ;
 wire \as2650.stack[8][1] ;
 wire \as2650.stack[8][2] ;
 wire \as2650.stack[8][3] ;
 wire \as2650.stack[8][4] ;
 wire \as2650.stack[8][5] ;
 wire \as2650.stack[8][6] ;
 wire \as2650.stack[8][7] ;
 wire \as2650.stack[8][8] ;
 wire \as2650.stack[8][9] ;
 wire \as2650.stack[9][0] ;
 wire \as2650.stack[9][10] ;
 wire \as2650.stack[9][11] ;
 wire \as2650.stack[9][12] ;
 wire \as2650.stack[9][13] ;
 wire \as2650.stack[9][14] ;
 wire \as2650.stack[9][15] ;
 wire \as2650.stack[9][1] ;
 wire \as2650.stack[9][2] ;
 wire \as2650.stack[9][3] ;
 wire \as2650.stack[9][4] ;
 wire \as2650.stack[9][5] ;
 wire \as2650.stack[9][6] ;
 wire \as2650.stack[9][7] ;
 wire \as2650.stack[9][8] ;
 wire \as2650.stack[9][9] ;
 wire \as2650.trap ;
 wire \as2650.warmup[0] ;
 wire \as2650.warmup[1] ;
 wire \as2650.wb_hidden_rom_enable ;
 wire clknet_0__01549_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf__01549_;
 wire clknet_1_1__leaf__01549_;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_136_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_leaf_146_wb_clk_i;
 wire clknet_leaf_147_wb_clk_i;
 wire clknet_leaf_148_wb_clk_i;
 wire clknet_leaf_149_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_150_wb_clk_i;
 wire clknet_leaf_151_wb_clk_i;
 wire clknet_leaf_152_wb_clk_i;
 wire clknet_leaf_153_wb_clk_i;
 wire clknet_leaf_154_wb_clk_i;
 wire clknet_leaf_155_wb_clk_i;
 wire clknet_leaf_157_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \wb_counter[0] ;
 wire \wb_counter[10] ;
 wire \wb_counter[11] ;
 wire \wb_counter[12] ;
 wire \wb_counter[13] ;
 wire \wb_counter[14] ;
 wire \wb_counter[15] ;
 wire \wb_counter[16] ;
 wire \wb_counter[17] ;
 wire \wb_counter[18] ;
 wire \wb_counter[19] ;
 wire \wb_counter[1] ;
 wire \wb_counter[20] ;
 wire \wb_counter[21] ;
 wire \wb_counter[22] ;
 wire \wb_counter[23] ;
 wire \wb_counter[24] ;
 wire \wb_counter[25] ;
 wire \wb_counter[26] ;
 wire \wb_counter[27] ;
 wire \wb_counter[28] ;
 wire \wb_counter[29] ;
 wire \wb_counter[2] ;
 wire \wb_counter[30] ;
 wire \wb_counter[31] ;
 wire \wb_counter[3] ;
 wire \wb_counter[4] ;
 wire \wb_counter[5] ;
 wire \wb_counter[6] ;
 wire \wb_counter[7] ;
 wire \wb_counter[8] ;
 wire \wb_counter[9] ;
 wire wb_debug_carry;
 wire wb_debug_cc;
 wire wb_feedback_delay;
 wire wb_io3_test;
 wire wb_reset_override;
 wire wb_reset_override_en;
 wire \web_behavior[0] ;
 wire \web_behavior[1] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05574__I (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05576__I (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__A1 (.I(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__A3 (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05581__A2 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05581__A3 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05582__I (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05583__A1 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__A1 (.I(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__A1 (.I(\as2650.indirect_target[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__A2 (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05588__I (.I(\as2650.PC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05589__A1 (.I(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__A2 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05594__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05594__A3 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05595__A1 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__A1 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05599__A4 (.I(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05600__A2 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05602__B2 (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__A1 (.I(\as2650.indirect_target[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__B2 (.I(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05604__A1 (.I(\as2650.indirect_target[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05604__B2 (.I(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__A1 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__A2 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__A3 (.I(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__A4 (.I(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__A1 (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05608__A1 (.I(\as2650.indirect_target[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05608__B2 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05610__B2 (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05611__A2 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05611__A3 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__B2 (.I(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__B1 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__B2 (.I(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__A2 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__A3 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05617__B1 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05619__A2 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05622__A2 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05623__A1 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05623__A2 (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05625__A2 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05625__B1 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05627__I (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__A1 (.I(\as2650.indirect_target[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__A2 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__B1 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__B2 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__I (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05632__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05635__A1 (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__A2 (.I(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__A2 (.I(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05638__I (.I(\as2650.instruction_args_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05640__A1 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05643__I (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05651__A1 (.I(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05652__I (.I(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05653__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05654__I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05656__A1 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05656__A2 (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05657__I (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05658__A1 (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05658__A2 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05659__I (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__A3 (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__A4 (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05663__A1 (.I(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__A1 (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__A2 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__A2 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05667__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05670__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05670__A3 (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05670__A4 (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05671__A1 (.I(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__A1 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__A2 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05674__A2 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05674__B (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05675__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05678__I (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__I (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__A2 (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05687__I (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05688__A2 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05688__A3 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05689__I (.I(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05693__I (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05695__I (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05697__A1 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__A1 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05700__A2 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05701__A1 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05702__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05703__S (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__I (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05713__A1 (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05715__I (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05716__I (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05717__I (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__A2 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__A2 (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__A3 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__B (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05721__I (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__A2 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05726__A1 (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__I (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A1 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A2 (.I(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__A1 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__A2 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__B1 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__B2 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__A1 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__I (.I(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05741__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__S (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__A1 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__A1 (.I(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05754__I (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__I (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I0 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I2 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I3 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__A1 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__A2 (.I(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__A4 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__A2 (.I(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__A2 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A1 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__I (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__A2 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05766__A2 (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__A1 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__A2 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A2 (.I(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__A2 (.I(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__A1 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__A2 (.I(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__A2 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__B2 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__I (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__S (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__I (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__A1 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__A1 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__I1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__I3 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__I (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__A2 (.I(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__A1 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__A2 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__B (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__S (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__I (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__A1 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__I0 (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__I1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__I2 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A2 (.I(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A4 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__I (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__I (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__I1 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__I3 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__B2 (.I(\as2650.PC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A1 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A2 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A3 (.I(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__A1 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A2 (.I(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__B1 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A2 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__A1 (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05836__I (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05837__S (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__A1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__A1 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__I (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__I0 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__I2 (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__I3 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__A4 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05854__A1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__A1 (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A1 (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A1 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__I (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I0 (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I2 (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I3 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__S0 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__S1 (.I(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__A1 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__A2 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__A1 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__A2 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__B (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A1 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A2 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A3 (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__A1 (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__S (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__I (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__A1 (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__A1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__A1 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__I (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I0 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I1 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I2 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I3 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__S0 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__A4 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A1 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A2 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__B (.I(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A1 (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__B1 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__B2 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05906__S (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__I (.I(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__A1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__A1 (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__I (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__I0 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__I1 (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__I3 (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__A2 (.I(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A1 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A2 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A2 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A3 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__I0 (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__I1 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__I2 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__I3 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A1 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A2 (.I(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A4 (.I(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__A2 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__B (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A1 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A2 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A2 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__B (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__A1 (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A2 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__B (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A2 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__A2 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__A2 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__A2 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A1 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A2 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A1 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A2 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A3 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A4 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__A1 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__B (.I(\as2650.instruction_args_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__A1 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A2 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__A1 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__A2 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__A1 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__A2 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A1 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__A1 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A1 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A2 (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__I (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__A1 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A1 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__A1 (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__A2 (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__I (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__I (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A1 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__I (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A1 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A1 (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A2 (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__I (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__A1 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__A3 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A2 (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__A4 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__A1 (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__A2 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A1 (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__I (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__A2 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__A1 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__A2 (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__A1 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__A1 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__A2 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__I (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__I (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__I (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__I (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__I (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__I (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__I (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__I (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__I (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__I (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__A2 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__I (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__A1 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__A4 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__I (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__A2 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__A2 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__B1 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__B2 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A1 (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__A2 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__B1 (.I(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__B2 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__C1 (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A1 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A2 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A2 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A3 (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__A2 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__A2 (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__A1 (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A1 (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A2 (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__A2 (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A2 (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A1 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A2 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A3 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A4 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__I (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__I (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__I (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A3 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A3 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A4 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A2 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__B (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__A1 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__A4 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__I (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__I (.I(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A2 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A3 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__A1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A1 (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A1 (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A2 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A2 (.I(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__I (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__I (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__I (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A1 (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__A1 (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__A2 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__A2 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__A1 (.I(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A1 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A2 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A2 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__I (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06189__A2 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A2 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__I (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A1 (.I(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A2 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__A1 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A2 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A2 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A3 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__I (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A2 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A1 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__I (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__A1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A2 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A1 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A2 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A2 (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A1 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A2 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__I (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A2 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A2 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A2 (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A3 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__I (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__I (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__I (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A2 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A3 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__A2 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A1 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A2 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A1 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__I (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__I (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A1 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A1 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A2 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A3 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A3 (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A3 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__A1 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A3 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__I (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__I (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A3 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__I (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A1 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__B (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A1 (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__I (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__I (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__I (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__I (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__I (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__I (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__I (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__I (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A2 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__I (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__I (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__I (.I(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__A1 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A1 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__A1 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A1 (.I(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A3 (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__I (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__A2 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__I (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__I (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__I (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A2 (.I(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A1 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__A1 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__A3 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__A4 (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A1 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A2 (.I(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A1 (.I(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A2 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A3 (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__A1 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__I (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A2 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__I (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__A2 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__I (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__I (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__I (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A1 (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A2 (.I(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A1 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__B (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A2 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A2 (.I(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__I (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A2 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__I (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A2 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__B (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A1 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A1 (.I(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__B (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__I (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__I (.I(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__I (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A1 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A2 (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__I (.I(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__I (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I0 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I1 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I2 (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I3 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__S0 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__S1 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__I (.I(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__I (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__I (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__I (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__I1 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__I3 (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__I (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06392__I1 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06392__I3 (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A1 (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A2 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A1 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A2 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A1 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A2 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__I (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__I1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__I3 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__I (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__I (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__A1 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A1 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__A1 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A1 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__B1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A1 (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A1 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A1 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I0 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I1 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I2 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I3 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A1 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A1 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A1 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__B1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A2 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__I (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__B1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__I (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A2 (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__A2 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A2 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A1 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A3 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A4 (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A2 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__A2 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__A1 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__B1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A3 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__B (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A1 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A2 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__I (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A2 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__I (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__A3 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__A4 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A3 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A4 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__I (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__A1 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__B (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__C (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A1 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A3 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06480__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A1 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A2 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__I (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A1 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__B2 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__C (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__A2 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__I (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__I (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A2 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A3 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__B1 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A1 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__A1 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__A2 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__I (.I(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A3 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A1 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A2 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A3 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__I (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__I (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A2 (.I(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A3 (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__I (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__B1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__B2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__I (.I(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__B (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__C (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A2 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A3 (.I(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__B (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__C (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A2 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__B (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__A1 (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__A2 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__B (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__I (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__C (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__I (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__I (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__I (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__I (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__I (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__I (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A3 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__I (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A1 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A2 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A2 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A2 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__A2 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A3 (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A1 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__B (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A1 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A2 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A3 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A1 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__I (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__I (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A2 (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__I (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__I (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A2 (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__I (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__I (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A1 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A3 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A2 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__B (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A1 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__C (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A1 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A4 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A1 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A2 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A2 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A1 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A2 (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__B1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__B2 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A1 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A2 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__I (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__A2 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__I (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__I (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__I (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A1 (.I(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A2 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__B1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__C (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A2 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__I (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__A1 (.I(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__A2 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A2 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__B1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__I (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__I (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__I (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__I (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__I (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__I (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A1 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A3 (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A2 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A3 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__I (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__I (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A1 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A4 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A2 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__A1 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__I (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A1 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A2 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A2 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A1 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__I (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__A1 (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A1 (.I(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A2 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A1 (.I(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A2 (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__A2 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__A1 (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__I (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A1 (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__A2 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A2 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A2 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A1 (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A2 (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A1 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A1 (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A2 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__I (.I(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__A2 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A2 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A1 (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__I (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__A1 (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A2 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A1 (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__A1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__I (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__I (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A2 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A2 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__A2 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A1 (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__I (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__A1 (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__I (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__I (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__A1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__A2 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A2 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A1 (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A1 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__I (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__A1 (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A2 (.I(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A2 (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A2 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__I (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A2 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__I (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A2 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__A2 (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A2 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A2 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__A1 (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__B1 (.I(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__B (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__I (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__I (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__I (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__I (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A1 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A2 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__I (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__I (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__I (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A2 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A3 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__I (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__I (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__A1 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__I (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A1 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__B (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__A2 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__I (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__I (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__I (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__I (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__I (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A2 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__I (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__I (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A1 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__B (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__I (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A2 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A1 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A1 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__I (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__I (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__I (.I(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__I (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A1 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__B (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A2 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__I (.I(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__I (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__C (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A1 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A2 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__I (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__I (.I(\as2650.PC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__I (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__I (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A1 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A2 (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A1 (.I(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A1 (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A1 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A2 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__I (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__I (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__I (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A1 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__C (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__I (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A2 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__I (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__I (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__C (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__I (.I(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__A1 (.I(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__I (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__I (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__I (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I (.I(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__A1 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__I (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__I (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__I (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__B (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A1 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__I (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__I (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__I (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A1 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__I (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A1 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__I (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__A2 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__I (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__I (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A1 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A1 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A2 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__I (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__I (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A1 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__I (.I(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__A1 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__A1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A2 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A2 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A2 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__I (.I(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A2 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__I (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A1 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A2 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A2 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__I (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__I (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A1 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A1 (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A2 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__I (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__I (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A1 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A1 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A2 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__I (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__I (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A1 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A1 (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A2 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__A1 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A1 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A2 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__I (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07056__I (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__A1 (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__A2 (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__I (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__I (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__I (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__I (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__I (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__I (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__I (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__I (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__I (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A1 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A1 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A1 (.I(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__I (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__I (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__I (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A1 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A2 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A3 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__I (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A3 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A4 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__I (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__B (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A1 (.I(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A2 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__I (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__I0 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__I1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__I0 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__I1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__I0 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__I1 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__I0 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__I1 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__I (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__I0 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__I1 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__I0 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__I1 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__I0 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__I1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__I0 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__I1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__I (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__I0 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__I1 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__I0 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__I1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__I1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__I0 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__I1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__I (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__I0 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__I1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__I0 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__I1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__I0 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__I1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__I0 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__I1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__I0 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__I1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__I0 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__I1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__I0 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__I1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__I0 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__I1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__I0 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__I1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__I0 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__I1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__I0 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__I1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__I0 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__I1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__I0 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__I1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__I0 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__I1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__I0 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__I1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__I0 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__I1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__I0 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__I1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__S (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__I0 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__I1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__S (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__I0 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__I1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__S (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__I0 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__I1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__S (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__I (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__I (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A1 (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A2 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__A2 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__I0 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__I1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__S (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__I0 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__I1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__S (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__I0 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__I1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__S (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__I (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A2 (.I(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__I (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A1 (.I(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A2 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A3 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__I (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__I (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__I (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A1 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A2 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__B (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A2 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__I (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__I (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A1 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A1 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__B (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A1 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A2 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__B (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A1 (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__I (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__I (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A2 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__A2 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__B (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A2 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__I (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__I (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A2 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A2 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__I (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A1 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A2 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A1 (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A2 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__B (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__I (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A2 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__I (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__I (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__A1 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A1 (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A2 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__B (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__A1 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__A2 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__I (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A2 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__A1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__A2 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__I (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__A2 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__I (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A3 (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__B (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__I (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A2 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__I (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__B (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__I (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__A1 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__B (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__B (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__I (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__I (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__I (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__A2 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__I (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A2 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A2 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__I (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__I (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A1 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A2 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A3 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__B1 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__B (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__C (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__I (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A2 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__B (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__B (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__I (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A2 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__B (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__I (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__B (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A2 (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A2 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__B (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__B (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__B (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A2 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__C (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__B (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__B (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A2 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A2 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__B1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A2 (.I(\wb_counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__B (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__C (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__B2 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__I (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__I (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__B1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__I (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__B1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A1 (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__B1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A1 (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__B1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A1 (.I(net287));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__B (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A2 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__B1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A1 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A2 (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__B (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A1 (.I(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__B1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__B2 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__C (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A1 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A1 (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A2 (.I(net427));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A1 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A2 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A1 (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A2 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A1 (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__C (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__I (.I(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__C (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__B (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__B (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__B (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__C (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__B (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__I (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__I (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__B (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__B (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__B (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__B (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__B (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__B (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__I (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__I (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__I (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__I (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__I (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A1 (.I(\wb_counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A2 (.I(\wb_counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__I (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__A1 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A1 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__I (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__A1 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A1 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A1 (.I(net392));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A2 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A1 (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A2 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__A2 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__B (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__A1 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__A2 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__I (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A1 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A2 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A1 (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A2 (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__B (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A1 (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A2 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A1 (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A2 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A2 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__A1 (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__A2 (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__B (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A1 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__I (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A2 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__I (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__I (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A2 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A2 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A3 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A2 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__I (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A2 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A3 (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__A1 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__I (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__B1 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A2 (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__I (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__I (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__I (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__I (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__I (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A1 (.I(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__C (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__I (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__I (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__I (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__I (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__I (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__I (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__I (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__C (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__B1 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__I (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__I (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__I (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__C (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__I (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__I (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__B1 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__I (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__I (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__I (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__C (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A1 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__I (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__I (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__I (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__I (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__S (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__I (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A1 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A3 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__B2 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__C1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__C2 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A2 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__I (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__I (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__I (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__I (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__I (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A2 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__I (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A1 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A3 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A2 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A1 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__I (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A1 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A2 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__I (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__B1 (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__B2 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__C (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A1 (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A2 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__I (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__I (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__B1 (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__B2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__C (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__I (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__I (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__I (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A1 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A2 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__I (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__I (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__B1 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__B2 (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__B (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__I (.I(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__I (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__B1 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__B2 (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__I (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__B (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__I (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__I (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__I (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__B1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__B2 (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__C (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__B1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__B2 (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__C (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__I (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A2 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A3 (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__I (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__I (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__I (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A2 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__I (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__I (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__I (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A2 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__B (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__B2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A2 (.I(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__I (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__I (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__I (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__I (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__I (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__C (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A2 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A2 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A3 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A4 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__I (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A2 (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A1 (.I(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A2 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__I (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__I (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__I (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__I (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A3 (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__I (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A1 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A2 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__B2 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A1 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__B2 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__C (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__C (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__I (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A1 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A2 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__I (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A1 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A1 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__I (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__B2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__I (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A1 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A2 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__I (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__A1 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__A2 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__B1 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A1 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__C (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__I (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A1 (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A2 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__I (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A2 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A2 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__A1 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__I (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A1 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__I (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__I (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__I (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A1 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A2 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__I (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__I (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__B2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__I (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A1 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A1 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__B2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A2 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__I (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__B1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__C (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__I (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__I (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A1 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A1 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__B1 (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A1 (.I(\as2650.indirect_target[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__B2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__I (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A1 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(\as2650.indirect_target[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A1 (.I(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A2 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__B (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__I (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__I (.I(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__I (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__I (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A1 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A2 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A2 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A2 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A2 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__I (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__I (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__I (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A1 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__B (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__B2 (.I(\as2650.indirect_target[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A1 (.I(\as2650.indirect_target[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A2 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__B (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__B (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__I (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__I (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A1 (.I(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__B (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__B2 (.I(\as2650.indirect_target[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A1 (.I(\as2650.indirect_target[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A2 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__B (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__B (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__I (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A1 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A2 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__B (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A1 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__B2 (.I(\as2650.indirect_target[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A1 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A2 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__B1 (.I(\as2650.indirect_target[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__B2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A1 (.I(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__B (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__I (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A1 (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__B1 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A1 (.I(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__I (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A1 (.I(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__B2 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__I (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A1 (.I(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A1 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A1 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A1 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A1 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A2 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__B2 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__A2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A1 (.I(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A1 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A2 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A3 (.I(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A4 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__I (.I(\as2650.instruction_args_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__I (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__B (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A1 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__A2 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__B1 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A1 (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A2 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A3 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A4 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__I (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A2 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A2 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__B1 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__B (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A1 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__B (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A1 (.I(\as2650.indirect_target[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__B2 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__C (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__A1 (.I(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__B (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A1 (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__I (.I(\as2650.instruction_args_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A2 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__C (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A1 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A3 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__I (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A4 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__B (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A3 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A1 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A2 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A1 (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__A1 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__I (.I(\as2650.instruction_args_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A3 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__B (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A1 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A2 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__B1 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A1 (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A2 (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A2 (.I(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A1 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__I (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__A2 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A1 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A2 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A2 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A1 (.I(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A1 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__I (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__B2 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__C (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__I (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A1 (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__B (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A1 (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__A1 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__A2 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__B1 (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A2 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__I (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A1 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__B1 (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A1 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__B2 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__I (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__B2 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A1 (.I(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A1 (.I(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__B2 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__I (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__I (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__B2 (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__B2 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A1 (.I(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A1 (.I(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__I (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A1 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__B2 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A1 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A1 (.I(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__I (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__I (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A2 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__B1 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__B1 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__I (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A2 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__B (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__I (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__I (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__B1 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A2 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__B (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__B2 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A3 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__B (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__I (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__B2 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__I (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A2 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__I (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__I (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__B2 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A2 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__I (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__B2 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A1 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A3 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A2 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__B2 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A1 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A3 (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__B1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__B2 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A1 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__I (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A3 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__I (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__B (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A1 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A2 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A3 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A1 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A3 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A1 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A2 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__C (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__I (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A1 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__A1 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A1 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A2 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__A1 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A1 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A2 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A3 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A1 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A2 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A2 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A1 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A2 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A1 (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A2 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A1 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A1 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A2 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A2 (.I(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A1 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__I (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__B2 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__C (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__I (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__I (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__B (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__I (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__B1 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__C (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__C (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__C (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__B1 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__I (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__C (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__S (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__B1 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__B (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A2 (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__B (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A1 (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__I (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__I (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__C (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__C (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__I (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__I (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__B1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__C (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__B1 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__I (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A1 (.I(\as2650.stack[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A2 (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__B1 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__C (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__S (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A1 (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__B1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A1 (.I(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A2 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__B (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A2 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A3 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__A1 (.I(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__A2 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__C (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A1 (.I(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__B (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A1 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__C (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__B (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__I (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A3 (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A4 (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A2 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__I (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__B (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A1 (.I(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__I (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__I (.I(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__B (.I(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__B (.I(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A1 (.I(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__B (.I(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A1 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__I (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__A1 (.I(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__B (.I(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A1 (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A2 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__I (.I(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__B (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A2 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__B (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A2 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__B (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A1 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A2 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A1 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__I (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A1 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A2 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__B (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A2 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__I (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__B2 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A2 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__B2 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__I (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__C (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__B2 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A2 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__B1 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__I (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__C (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__S (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A2 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A3 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__B (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__I (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A2 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A3 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__B (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A2 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__I (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__I (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A2 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__B2 (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__I (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__I (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A1 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__I (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__I (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__I (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A2 (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__B1 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__I (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__I (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__B1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__C (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__I (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__B1 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A2 (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__B1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__C (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__B1 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__B1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__C (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A2 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__B1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A2 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__B1 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__C (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__I (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__S (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A2 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A3 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__B1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__B2 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__A2 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__B (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A2 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A1 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A2 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A1 (.I(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__A2 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__I (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A2 (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__B1 (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__C (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__B1 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A2 (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__B1 (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__C (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__C (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__B1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__B1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__C (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A1 (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__I0 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__S (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__B1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A1 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A2 (.I(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A2 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__B (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__A2 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__B1 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A2 (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__B1 (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__C (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A2 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__B1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__C (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A2 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A2 (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__B1 (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__C (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__B1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__B1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__C (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__S (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A2 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A2 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A2 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__B2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__B1 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__B2 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__C (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__B1 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__C (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__B1 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__B2 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__B2 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__C (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__B1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A2 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__B1 (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__C (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__S (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__B1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__B2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A1 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__B1 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__B2 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__C (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A2 (.I(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A2 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__B1 (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__B2 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__C (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__C (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__B1 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__B1 (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__B2 (.I(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__C (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A2 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__B1 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A2 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__C (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A1 (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__S (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A2 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__B2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__C (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A2 (.I(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A1 (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A2 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__B (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A3 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A1 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A2 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A1 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__I (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__B2 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__C (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A1 (.I(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__B1 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__B2 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__C (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__I (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A2 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__B1 (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__C (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A1 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__S (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A1 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__B1 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__B2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A2 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__A1 (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__B (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A1 (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A2 (.I(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__I (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__B1 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__B2 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__B2 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__B1 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__C (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__B1 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__B2 (.I(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__B1 (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__B2 (.I(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__B1 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__B2 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__C (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__S (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A2 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__B2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__C (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A1 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A1 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__B (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A3 (.I(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A2 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A3 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__I (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__I (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A2 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__B1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__C (.I(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__I (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A1 (.I(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__B1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__B2 (.I(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__C (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A2 (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__B1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__C (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A2 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__B1 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__B1 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__C (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A1 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__S (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__B1 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__C (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A2 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__B2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A2 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__B1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A2 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__B1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__C (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__B1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__C (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__B2 (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A1 (.I(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__B1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__B2 (.I(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__C (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__B2 (.I(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__B1 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__B2 (.I(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__C (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__S (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__B1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A2 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__B1 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__C (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__B2 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__C (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A1 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A2 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A2 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A2 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A2 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__B2 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__I (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__B1 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A2 (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__B1 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__C (.I(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__B1 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__C (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__B2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__B1 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A2 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__B1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__C (.I(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A2 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__B1 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A2 (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__B1 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__C (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__S (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__B1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A1 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A2 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__B (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__I (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__C (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A2 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__B (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A2 (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__B1 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__B1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__C (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__B1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__C (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__B2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__B2 (.I(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__C (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__B1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__B2 (.I(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__B2 (.I(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__C (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__S (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__B1 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A1 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A2 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A2 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__B2 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A2 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A2 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__B (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A2 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A3 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__B1 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A2 (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__B1 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__C (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__B1 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A2 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__B1 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__C (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__B1 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__B1 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__C (.I(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A2 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__B1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A2 (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__B1 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__C (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__S (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__B1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A2 (.I(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__B (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__C (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__C (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__C (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A2 (.I(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__I (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A1 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A2 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A2 (.I(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A2 (.I(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A1 (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A2 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A2 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A2 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A1 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A2 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A2 (.I(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A1 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A1 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A1 (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A1 (.I(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A2 (.I(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A2 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__I0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__I0 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__I1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__S (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A2 (.I(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__I (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A2 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A1 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A2 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A2 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A2 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A1 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__I (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__I (.I(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A1 (.I(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__B (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__I (.I(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__I (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A1 (.I(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__I0 (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__B (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A2 (.I(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__I (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A2 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__C (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__I (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A2 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__B (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__C (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A1 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__B1 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__I (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A2 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__I (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__I (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__I (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A1 (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A2 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__I (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A1 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A3 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__I (.I(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A2 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A3 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__I (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__B (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A2 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__B (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__B (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A1 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A3 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A2 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A3 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__I (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__B2 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A1 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__B (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A1 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__C (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__I (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__I (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A2 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__B2 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__B (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A1 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A2 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__B2 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A1 (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A2 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A2 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A2 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__I (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A3 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A2 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__I (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A3 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__I (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__I (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A1 (.I(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__B (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__C (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A1 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__B1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__I (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A1 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A1 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__C (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A1 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A1 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A3 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A2 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__B (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A1 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A3 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A2 (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__B2 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A1 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A2 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A1 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__B (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__B2 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__I (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__I (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A1 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A1 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A1 (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A2 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A2 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__B (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A2 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A1 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__C (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A3 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A2 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A2 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A1 (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__I (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__I (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__I (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__B2 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A1 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__B1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__B2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__C (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A1 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A2 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A2 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__A2 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A1 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A2 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__A2 (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A1 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A2 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A1 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__B1 (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__B2 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A2 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A4 (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A1 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A2 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__A1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A2 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__B2 (.I(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A1 (.I(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A1 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A2 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A2 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A1 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A2 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A2 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A1 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A2 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A1 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A2 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A2 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A2 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A2 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__B1 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__B2 (.I(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A3 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A4 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A2 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A2 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A2 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A2 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A1 (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09328__A1 (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A2 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__B2 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__A2 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A1 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A2 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A2 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A4 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A2 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A1 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__B2 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A1 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A2 (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A1 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A1 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A1 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A2 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A1 (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A2 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__B (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__C (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A2 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A2 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A2 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A3 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A2 (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A1 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A2 (.I(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A2 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A1 (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A1 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__I (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A1 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A2 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A3 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A1 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A2 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A3 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A3 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__B2 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A1 (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__A1 (.I(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__C (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A2 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__B1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__B1 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__C (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__C (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A2 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__B1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__C (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A2 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__B1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A1 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A2 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A4 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A1 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__B1 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__C (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A1 (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__B1 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__C (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__B1 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__B2 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A2 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__B1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__A1 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__B1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__B2 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__B1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__B2 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A2 (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A2 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A1 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A1 (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A1 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A2 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__B2 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A2 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A1 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A1 (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A2 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__B (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__I (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__I (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A2 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A3 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A4 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A1 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A2 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__B (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A1 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A2 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A2 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A3 (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A2 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A2 (.I(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A3 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A2 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A3 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A4 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A2 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A2 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A2 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__B (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__C (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A2 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__A1 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__I0 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__I1 (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A1 (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A2 (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A2 (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A1 (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__A1 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A2 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A1 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__B2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A2 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__B2 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A1 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A2 (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A3 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A2 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A2 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__B1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__B2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09655__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09655__A2 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A1 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__B1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__C1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__C2 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A2 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__B (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__C (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__B1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__B2 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A1 (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A1 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A2 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A3 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A2 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__B1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__B2 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A2 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__B1 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__B2 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__I (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A2 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B2 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A2 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__B1 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__B2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__B1 (.I(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__I (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A2 (.I(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__B (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A1 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A2 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__B (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__B (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A2 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__I (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A1 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A2 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__B (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A1 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A2 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A3 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A4 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A3 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A3 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A1 (.I(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A2 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__C (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I0 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I3 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__I0 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__I1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__I2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__I1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__I2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__S1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__I0 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__I2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__I1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__I2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__I0 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__I1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__I2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__S1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A3 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A4 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A2 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A3 (.I(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__I2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A1 (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A2 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__B (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A3 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A1 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__B1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__B2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__B (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__C (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A1 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A3 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A2 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A1 (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A2 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__B2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__B (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__B (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A2 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__B (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__I (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__B (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__C (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A2 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A3 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__C (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A2 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__I (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A2 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__A1 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A2 (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__B (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A1 (.I(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A1 (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A1 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A1 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A1 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A2 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A2 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A3 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__B2 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A2 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A1 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A1 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A2 (.I(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__I0 (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A1 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A1 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A1 (.I(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A3 (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__B2 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__A1 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__A3 (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__A1 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__B (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__B2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A1 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A1 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__B2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__C (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A2 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A3 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A1 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__B2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__I (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__C (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A2 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A3 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A1 (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__B (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A1 (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__I (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__I0 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__I0 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__I0 (.I(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__I0 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__I0 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__S (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__I0 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__S (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__I (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A1 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__I (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__I (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A1 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A1 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__I (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A2 (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A2 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A3 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__B2 (.I(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A1 (.I(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__I (.I(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A2 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A2 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A2 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A2 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A2 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__A2 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__A2 (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A2 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__I (.I(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A2 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A2 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A2 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A2 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A2 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A2 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A2 (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A2 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__A2 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A1 (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A2 (.I(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__I (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A1 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__I (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__A1 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__I (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A1 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A1 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A2 (.I(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__B (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A2 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__B (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__B (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A1 (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A2 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__A1 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__A1 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__B (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A2 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A1 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__A1 (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__B (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A2 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__I (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__I (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A2 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A2 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A2 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A2 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A2 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A2 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A2 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A2 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__I (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__I (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__I (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__I (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A1 (.I(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__A1 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A1 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__I (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__I (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A2 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A2 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A2 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A2 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__I (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__I (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__A1 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__I (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A1 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__I (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__I (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__I (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A1 (.I(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__I (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A1 (.I(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__I (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__I (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__I (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__I (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__I (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__I (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A2 (.I(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A2 (.I(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__I (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A2 (.I(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A2 (.I(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A2 (.I(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A2 (.I(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__I (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A2 (.I(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__A2 (.I(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__I (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__I (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A1 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__I (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__I (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__I (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__I (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__I (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__I (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A2 (.I(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__B (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A2 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A2 (.I(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A3 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A1 (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A2 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A1 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A2 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A1 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__I (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A3 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A1 (.I(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A3 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A2 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A3 (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A4 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__A1 (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A2 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A3 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A3 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__A2 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A1 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A1 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A2 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__B1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__B2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__C (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A2 (.I(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__B (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A1 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A2 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__A1 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__I (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__I (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__I (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A2 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__I (.I(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A2 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__I (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__B (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A2 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__B2 (.I(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__I (.I(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__C (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__I (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A2 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A2 (.I(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__C (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__I (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A2 (.I(\as2650.instruction_args_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__B (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A1 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A2 (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__I (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A3 (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__I (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__A2 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__I (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__I (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__I (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A2 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A2 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__A1 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__I (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A1 (.I(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A1 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__C (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A2 (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__B2 (.I(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__I (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__I (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__I (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__I (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A2 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A3 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__B (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__B2 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A2 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A3 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A4 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__A1 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__I (.I(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A1 (.I(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A2 (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A3 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__I (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A1 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__I (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__A1 (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__C (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A1 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A2 (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__C (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A1 (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A1 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A1 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__B1 (.I(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__C1 (.I(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__I (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A2 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__I (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__I (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__B (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A1 (.I(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__B2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__I (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__I (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__I (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A1 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__I (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A2 (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__B2 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__C (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__C (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__A1 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A1 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A1 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__B1 (.I(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__C1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__I (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__I (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__B (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__B2 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A2 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__A1 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A1 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A2 (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__C (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__C (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A1 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A1 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__B1 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__C1 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__I (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A1 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__B (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__B2 (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A2 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A3 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__C (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A1 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A2 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A1 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__A1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__B1 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__C (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__A1 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__A2 (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__B (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A1 (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A1 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A1 (.I(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A1 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__B1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__C1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__I (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A1 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__B (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__B2 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A1 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A1 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__B (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__I (.I(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A1 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__C (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A2 (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A2 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A1 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A1 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__I (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__B1 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__C1 (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__B (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A1 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__B2 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A2 (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__B (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A1 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__B2 (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__C (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__C (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A3 (.I(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A1 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__A1 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A1 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__A1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__B1 (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__C1 (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__B (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__B2 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__A2 (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__B (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A1 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A1 (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A1 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__B (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A2 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A2 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__C (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A2 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__B (.I(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A1 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__B1 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__C1 (.I(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__I (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__I (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__I (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__A1 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__I (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__I (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__I (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__I (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__I (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__I (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A2 (.I(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A2 (.I(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A2 (.I(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A2 (.I(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A1 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A2 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A2 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A2 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A2 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A2 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A2 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__A2 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A2 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__I (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__I (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__A1 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__I (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__A1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A1 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__I (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__I (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__I (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A2 (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A2 (.I(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__I (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A2 (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__A2 (.I(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A2 (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A2 (.I(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__I (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A2 (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A1 (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A2 (.I(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__I (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__I (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__I (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__I (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A1 (.I(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__I (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__I (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__I (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A2 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A2 (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__I (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A2 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A2 (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__A2 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__A2 (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__I (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A1 (.I(\as2650.stack[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A2 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__A2 (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__I (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__I (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A1 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__A1 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__I (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__I (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__A1 (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__I (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__I (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A1 (.I(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__I (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__I (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A2 (.I(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A2 (.I(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__A2 (.I(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A2 (.I(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__I (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A1 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A2 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A1 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__A1 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__A2 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A1 (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__B2 (.I(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A1 (.I(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__B2 (.I(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A1 (.I(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__B2 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A1 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__B2 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__B2 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A1 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__B2 (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__A1 (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__B2 (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A1 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__B2 (.I(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__I (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A2 (.I(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__B (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A1 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__I (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__I (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A2 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__I (.I(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__I (.I(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__I (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__I (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__I (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A1 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__I (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__I (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__I (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__I (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__I (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__A1 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__I (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__I (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__I (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__A1 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__A2 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A2 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A1 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A2 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A2 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__I (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__I (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A1 (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__I (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__I (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A1 (.I(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A1 (.I(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__I (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__I (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A2 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A2 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A2 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A2 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A2 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A2 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A2 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A2 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A3 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A2 (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A1 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A1 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__A1 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__A1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A1 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__A1 (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A1 (.I(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A2 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A2 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__A2 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__A2 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A2 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A1 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A2 (.I(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A1 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A2 (.I(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A1 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A2 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A2 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__I (.I(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__I (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__I1 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A2 (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A2 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__A1 (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__A2 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A1 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A2 (.I(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A3 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__I (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__I (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A3 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__A2 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__A2 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__I (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A1 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__I1 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__A2 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A2 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__A1 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A1 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A2 (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A1 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A2 (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A1 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A1 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A2 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__B1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A1 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__A2 (.I(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A1 (.I(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A2 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__B1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A1 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A1 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A3 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A1 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A1 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A2 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__B1 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A2 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A3 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A1 (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__A1 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A2 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A3 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A2 (.I(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A1 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A2 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__I (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A3 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A1 (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A2 (.I(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A2 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A3 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A2 (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A1 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A1 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A2 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A3 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__I (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A1 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__B1 (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A3 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A1 (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A3 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A1 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A3 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__B (.I(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A3 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A2 (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A1 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A1 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A2 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A1 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A2 (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A3 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A1 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A2 (.I(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A2 (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A1 (.I(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__I (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__I (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A2 (.I(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A2 (.I(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__I (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__A2 (.I(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A2 (.I(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__A2 (.I(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A2 (.I(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A2 (.I(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A2 (.I(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__I (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__I (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__I (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__I (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A1 (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__I (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A1 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__I (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__I (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__I (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A1 (.I(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__I (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A1 (.I(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__I (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__I (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__I (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__I (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A1 (.I(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__I (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__A3 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__I (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__A2 (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__I (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__A1 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__I (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__I (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A2 (.I(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A2 (.I(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A2 (.I(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__A2 (.I(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A2 (.I(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A2 (.I(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A2 (.I(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__A2 (.I(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__I (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__I (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__A1 (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A1 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A1 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__I (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__I (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A1 (.I(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A1 (.I(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A1 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__A1 (.I(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__A1 (.I(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__I (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__I (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__I (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__I (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__I (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__I (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A1 (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__A1 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__A1 (.I(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A1 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__I (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__I (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A1 (.I(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A1 (.I(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__A1 (.I(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A1 (.I(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__I (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__I (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__I (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__I (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A2 (.I(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A2 (.I(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A2 (.I(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__A2 (.I(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A2 (.I(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A2 (.I(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A2 (.I(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A2 (.I(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__I (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__I (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A1 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A1 (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A1 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__I (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__I (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A1 (.I(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A1 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A1 (.I(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A1 (.I(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__I (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__I (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__A2 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A2 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A2 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A2 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__CLK (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__D (.I(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__D (.I(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__D (.I(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__D (.I(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__D (.I(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__D (.I(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__D (.I(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__D (.I(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__D (.I(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__D (.I(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11581__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__CLK (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11649__CLK (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11650__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11652__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11855__I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11856__I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__I (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11858__I (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11859__I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11860__I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11861__I (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_136_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_137_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_140_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_142_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_146_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_147_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_148_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_149_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_150_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_151_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_152_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_153_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_154_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_155_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_157_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold100_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold101_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold102_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold103_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold104_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold105_I (.I(wbs_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold106_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold107_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold108_I (.I(wbs_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold109_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold110_I (.I(wbs_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold111_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold112_I (.I(wbs_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold113_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold114_I (.I(wbs_adr_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold115_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold116_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold117_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold118_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold119_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold120_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold121_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold14_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold18_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold22_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold28_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold33_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold37_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold42_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold44_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold46_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold48_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold50_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold52_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold54_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold56_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold58_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold60_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold66_I (.I(wbs_adr_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold67_I (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold82_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold83_I (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold84_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold85_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold86_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold88_I (.I(wbs_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold89_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold90_I (.I(wbs_adr_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold91_I (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold92_I (.I(wbs_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold93_I (.I(wbs_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold94_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold95_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold96_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold97_I (.I(wbs_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold98_I (.I(wbs_adr_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold99_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(bus_in_serial_ports[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(bus_in_serial_ports[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(bus_in_serial_ports[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(bus_in_serial_ports[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(bus_in_serial_ports[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(bus_in_serial_ports[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(bus_in_serial_ports[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(bus_in_sid[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(bus_in_sid[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(bus_in_sid[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(bus_in_gpios[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(bus_in_sid[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(bus_in_sid[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(bus_in_sid[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(bus_in_sid[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(bus_in_sid[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(bus_in_timers[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(bus_in_timers[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(bus_in_timers[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(bus_in_timers[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(bus_in_timers[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(bus_in_gpios[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(bus_in_timers[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(bus_in_timers[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(bus_in_timers[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(bus_in_gpios[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(irqs[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(irqs[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(irqs[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(irqs[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(irqs[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(irqs[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(irqs[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(bus_in_gpios[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(ram_bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(ram_bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(ram_bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(ram_bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(ram_bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(ram_bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(ram_bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(ram_bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(rom_bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(rom_bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(bus_in_gpios[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(rom_bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(rom_bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(rom_bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(rom_bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(rom_bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(rom_bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(bus_in_gpios[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_in_gpios[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(bus_in_gpios[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(bus_in_serial_ports[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap304_I (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output132_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output133_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output134_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output155_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output156_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output196_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output198_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output199_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output200_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output209_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output210_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output211_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output212_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output213_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output214_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output215_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output216_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output217_I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output218_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output219_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output220_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output221_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output223_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output224_I (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output225_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output226_I (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output227_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output230_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output231_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output234_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output236_I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output237_I (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output238_I (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output239_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output241_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output242_I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output243_I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output244_I (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output245_I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output246_I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output247_I (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output248_I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output249_I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output250_I (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output251_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output252_I (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output253_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output254_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output255_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output256_I (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output266_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output276_I (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output277_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output281_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output282_I (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output283_I (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output284_I (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output285_I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output286_I (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output287_I (.I(net287));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output288_I (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output289_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output290_I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output291_I (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output292_I (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output293_I (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer12_I (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer2_I (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer3_I (.I(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire298_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire299_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire300_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_627 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05574_ (.I(\as2650.cycle[9] ),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05575_ (.I(_00588_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05576_ (.I(_00589_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05577_ (.I(_00590_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05578_ (.I(\as2650.PC[7] ),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05579_ (.A1(\as2650.relative_cyc ),
    .A2(\as2650.indirect_cyc ),
    .A3(\as2650.cycle[9] ),
    .A4(\as2650.is_interrupt_cycle ),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05580_ (.I(_00593_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05581_ (.A1(\as2650.cycle[0] ),
    .A2(\as2650.cycle[4] ),
    .A3(\as2650.cycle[6] ),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05582_ (.I(_00595_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05583_ (.A1(_00594_),
    .A2(_00596_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05584_ (.A1(\as2650.relative_cyc ),
    .A2(\as2650.indirect_cyc ),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05585_ (.I(_00598_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05586_ (.A1(\as2650.indirect_target[7] ),
    .A2(_00599_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05587_ (.A1(_00592_),
    .A2(_00597_),
    .B(_00600_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05588_ (.I(\as2650.PC[3] ),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05589_ (.A1(\as2650.relative_cyc ),
    .A2(\as2650.indirect_cyc ),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05590_ (.I(\as2650.indirect_target[3] ),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _05591_ (.A1(_00602_),
    .A2(_00594_),
    .A3(_00596_),
    .B1(_00603_),
    .B2(_00604_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05592_ (.I(\as2650.PC[1] ),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05593_ (.I(\as2650.indirect_target[1] ),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _05594_ (.A1(_00606_),
    .A2(_00593_),
    .A3(_00595_),
    .B1(_00603_),
    .B2(_00607_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05595_ (.A1(\as2650.cycle[4] ),
    .A2(\as2650.indirect_target[0] ),
    .A3(_00598_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05596_ (.I(\as2650.PC[2] ),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05597_ (.I(\as2650.indirect_target[2] ),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _05598_ (.A1(_00610_),
    .A2(_00593_),
    .A3(_00596_),
    .B1(_00603_),
    .B2(_00611_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05599_ (.A1(_00605_),
    .A2(_00608_),
    .A3(_00609_),
    .A4(_00612_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05600_ (.A1(_00593_),
    .A2(_00595_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05601_ (.I(_00614_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05602_ (.A1(\as2650.indirect_target[4] ),
    .A2(_00599_),
    .B1(_00615_),
    .B2(\as2650.PC[4] ),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05603_ (.A1(\as2650.indirect_target[5] ),
    .A2(_00598_),
    .B1(_00614_),
    .B2(\as2650.PC[5] ),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05604_ (.A1(\as2650.indirect_target[6] ),
    .A2(_00599_),
    .B1(_00615_),
    .B2(\as2650.PC[6] ),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05605_ (.A1(_00613_),
    .A2(_00616_),
    .A3(_00617_),
    .A4(_00618_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05606_ (.A1(_00601_),
    .A2(_00619_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05607_ (.I(_00599_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05608_ (.A1(\as2650.indirect_target[8] ),
    .A2(_00621_),
    .B1(_00615_),
    .B2(\as2650.PC[8] ),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05609_ (.I(_00615_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05610_ (.A1(\as2650.indirect_target[9] ),
    .A2(_00621_),
    .B1(_00623_),
    .B2(\as2650.PC[9] ),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05611_ (.A1(_00620_),
    .A2(_00622_),
    .A3(_00624_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05612_ (.I(_00621_),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05613_ (.A1(\as2650.indirect_target[10] ),
    .A2(_00626_),
    .B1(_00623_),
    .B2(\as2650.PC[10] ),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05614_ (.I(_00623_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05615_ (.A1(\as2650.indirect_target[11] ),
    .A2(_00626_),
    .B1(_00628_),
    .B2(\as2650.PC[11] ),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05616_ (.A1(_00625_),
    .A2(_00627_),
    .A3(_00629_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05617_ (.A1(\as2650.indirect_target[12] ),
    .A2(_00626_),
    .B1(_00628_),
    .B2(\as2650.PC[12] ),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05618_ (.I(_00631_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05619_ (.A1(_00630_),
    .A2(_00632_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05620_ (.I(\as2650.page_reg[0] ),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05621_ (.I(_00626_),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05622_ (.A1(\as2650.indirect_target[13] ),
    .A2(_00635_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05623_ (.A1(_00634_),
    .A2(_00597_),
    .B(_00636_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05624_ (.A1(_00633_),
    .A2(_00637_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05625_ (.A1(\as2650.indirect_target[14] ),
    .A2(_00635_),
    .B1(_00628_),
    .B2(\as2650.page_reg[1] ),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05626_ (.A1(_00638_),
    .A2(_00639_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05627_ (.I(_00628_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05628_ (.A1(\as2650.indirect_target[15] ),
    .A2(_00635_),
    .B1(_00641_),
    .B2(\as2650.page_reg[2] ),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05629_ (.A1(_00640_),
    .A2(_00642_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05630_ (.I(\as2650.page_reg[2] ),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05631_ (.I(\as2650.indirect_cyc ),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05632_ (.A1(_00645_),
    .A2(\as2650.extend ),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05633_ (.I(_00646_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05634_ (.A1(\as2650.instruction_args_latch[15] ),
    .A2(_00647_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05635_ (.A1(_00644_),
    .A2(_00647_),
    .B(_00648_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05636_ (.A1(_00591_),
    .A2(_00649_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05637_ (.A1(_00591_),
    .A2(_00643_),
    .B(_00650_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05638_ (.I(\as2650.instruction_args_latch[14] ),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05639_ (.A1(\as2650.page_reg[1] ),
    .A2(_00646_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05640_ (.A1(_00652_),
    .A2(_00647_),
    .B(_00653_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05641_ (.A1(_00638_),
    .A2(_00639_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05642_ (.I0(_00654_),
    .I1(_00655_),
    .S(_00591_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05643_ (.I(\as2650.cycle[9] ),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05644_ (.A1(\as2650.indexed_cyc[1] ),
    .A2(\as2650.indexed_cyc[0] ),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05645_ (.I(_00658_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05646_ (.A1(_00657_),
    .A2(_00659_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05647_ (.I(_00660_),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05648_ (.I(_00661_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05649_ (.I(\as2650.cycle[0] ),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05650_ (.I(_00663_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05651_ (.A1(\as2650.wb_hidden_rom_enable ),
    .A2(\as2650.cpu_hidden_rom_enable ),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05652_ (.I(_00665_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _05653_ (.A1(net59),
    .A2(_00666_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05654_ (.I(net239),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05655_ (.I(_00668_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _05656_ (.A1(net227),
    .A2(net226),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05657_ (.I(_00670_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _05658_ (.A1(net225),
    .A2(net224),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05659_ (.I(_00672_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05660_ (.I(net39),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05661_ (.A1(_00669_),
    .A2(_00671_),
    .A3(_00673_),
    .B(_00674_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _05662_ (.A1(_00668_),
    .A2(net51),
    .A3(_00670_),
    .A4(_00672_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _05663_ (.A1(_00665_),
    .A2(_00675_),
    .A3(_00676_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05664_ (.A1(_00667_),
    .A2(_00677_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05665_ (.A1(\as2650.insin[1] ),
    .A2(_00663_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05666_ (.A1(_00664_),
    .A2(_00678_),
    .B(_00679_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _05667_ (.A1(net58),
    .A2(_00666_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05668_ (.I(net38),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05669_ (.A1(_00669_),
    .A2(_00671_),
    .A3(_00673_),
    .B(_00682_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _05670_ (.A1(_00669_),
    .A2(net50),
    .A3(_00670_),
    .A4(_00672_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _05671_ (.A1(_00665_),
    .A2(_00683_),
    .A3(_00684_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05672_ (.A1(_00681_),
    .A2(_00685_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05673_ (.A1(\as2650.insin[0] ),
    .A2(_00663_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05674_ (.A1(_00663_),
    .A2(_00686_),
    .B(_00687_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05675_ (.I(\as2650.debug_psl[4] ),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05676_ (.I(_00689_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05677_ (.I(_00690_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05678_ (.I(_00691_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05679_ (.I(_00692_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05680_ (.I(_00693_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05681_ (.I(\as2650.regs[3][7] ),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05682_ (.A1(_00694_),
    .A2(\as2650.regs[7][7] ),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05683_ (.A1(_00694_),
    .A2(_00695_),
    .B(_00696_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05684_ (.A1(_00688_),
    .A2(_00697_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05685_ (.I(\as2650.cycle[0] ),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05686_ (.I(_00699_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05687_ (.I(_00687_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05688_ (.A1(_00700_),
    .A2(_00681_),
    .A3(_00685_),
    .B(_00701_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05689_ (.I(_00702_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05690_ (.I(_00703_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05691_ (.I(_00704_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05692_ (.I(_00705_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05693_ (.I(_00691_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05694_ (.I(_00707_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05695_ (.I(_00708_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05696_ (.I(\as2650.regs[2][7] ),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05697_ (.A1(_00709_),
    .A2(\as2650.regs[6][7] ),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05698_ (.A1(_00709_),
    .A2(_00710_),
    .B(_00711_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05699_ (.I(_00712_),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05700_ (.A1(_00706_),
    .A2(net203),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05701_ (.A1(_00680_),
    .A2(_00698_),
    .A3(_00713_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05702_ (.I(\as2650.debug_psl[4] ),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05703_ (.I0(\as2650.regs[1][7] ),
    .I1(\as2650.regs[5][7] ),
    .S(_00715_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05704_ (.I(_00716_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05705_ (.I(_00717_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05706_ (.I(_00718_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05707_ (.I(_00719_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05708_ (.I(_00720_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _05709_ (.I(_00721_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05710_ (.I(_00690_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05711_ (.I(_00723_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05712_ (.I(\as2650.regs[0][7] ),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05713_ (.A1(_00691_),
    .A2(_00725_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05714_ (.A1(_00724_),
    .A2(\as2650.regs[4][7] ),
    .B(_00726_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05715_ (.I(_00727_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05716_ (.I(_00728_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05717_ (.I(_00729_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05718_ (.A1(_00705_),
    .A2(_00730_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05719_ (.I(_00679_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05720_ (.A1(_00699_),
    .A2(_00667_),
    .A3(_00677_),
    .B(_00732_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05721_ (.I(net345),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05722_ (.I(_00734_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05723_ (.I(_00735_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05724_ (.A1(_00706_),
    .A2(_00722_),
    .B(_00731_),
    .C(_00736_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05725_ (.A1(_00714_),
    .A2(_00737_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05726_ (.A1(_00601_),
    .A2(net430),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05727_ (.I(_00620_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05728_ (.A1(_00590_),
    .A2(_00740_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05729_ (.I(_00588_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05730_ (.I(_00742_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05731_ (.I(_00743_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05732_ (.I(_00744_),
    .Z(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05733_ (.A1(_00745_),
    .A2(\as2650.instruction_args_latch[7] ),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05734_ (.A1(_00662_),
    .A2(_00738_),
    .B1(_00739_),
    .B2(_00741_),
    .C(_00746_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05735_ (.I(_00743_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05736_ (.I(_00659_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05737_ (.I(\as2650.regs[3][6] ),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05738_ (.A1(_00693_),
    .A2(\as2650.regs[7][6] ),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05739_ (.A1(_00709_),
    .A2(_00750_),
    .B(_00751_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05740_ (.I(_00752_),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05741_ (.I(\as2650.debug_psl[4] ),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05742_ (.I0(\as2650.regs[1][6] ),
    .I1(\as2650.regs[5][6] ),
    .S(_00753_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05743_ (.I(_00754_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05744_ (.I(_00755_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05745_ (.I(_00756_),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05746_ (.I(_00757_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05747_ (.I(\as2650.regs[2][6] ),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05748_ (.A1(_00709_),
    .A2(\as2650.regs[6][6] ),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05749_ (.A1(_00694_),
    .A2(_00759_),
    .B(_00760_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05750_ (.I(_00761_),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05751_ (.I(\as2650.regs[0][6] ),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05752_ (.A1(_00690_),
    .A2(_00762_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05753_ (.A1(_00691_),
    .A2(\as2650.regs[4][6] ),
    .B(_00763_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05754_ (.I(_00764_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05755_ (.I(_00765_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05756_ (.I(_00766_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05757_ (.I(_00704_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05758_ (.I0(net211),
    .I1(_00758_),
    .I2(net202),
    .I3(_00767_),
    .S0(_00735_),
    .S1(_00768_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05759_ (.A1(_00748_),
    .A2(\as2650.instruction_args_latch[6] ),
    .A3(_00749_),
    .A4(_00769_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05760_ (.A1(_00688_),
    .A2(_00752_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05761_ (.A1(_00705_),
    .A2(net202),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05762_ (.A1(_00680_),
    .A2(_00771_),
    .A3(_00772_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _05763_ (.I(_00758_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05764_ (.I(_00766_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05765_ (.A1(_00768_),
    .A2(_00775_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05766_ (.A1(_00705_),
    .A2(_00774_),
    .B(_00776_),
    .C(_00736_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05767_ (.A1(_00773_),
    .A2(_00777_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05768_ (.A1(_00613_),
    .A2(_00616_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05769_ (.A1(_00779_),
    .A2(_00617_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05770_ (.A1(_00780_),
    .A2(_00618_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05771_ (.A1(_00748_),
    .A2(\as2650.instruction_args_latch[6] ),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05772_ (.A1(_00661_),
    .A2(_00778_),
    .B1(_00781_),
    .B2(_00748_),
    .C(_00782_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05773_ (.A1(_00770_),
    .A2(_00783_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05774_ (.I(\as2650.regs[3][5] ),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05775_ (.A1(_00693_),
    .A2(\as2650.regs[7][5] ),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05776_ (.A1(_00693_),
    .A2(_00785_),
    .B(_00786_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05777_ (.I(_00787_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05778_ (.I(_00689_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05779_ (.I0(\as2650.regs[1][5] ),
    .I1(\as2650.regs[5][5] ),
    .S(_00789_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05780_ (.I(_00790_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05781_ (.I(_00791_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05782_ (.I(_00792_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05783_ (.I(_00793_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05784_ (.I(\as2650.regs[2][5] ),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05785_ (.I(_00724_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05786_ (.A1(_00796_),
    .A2(\as2650.regs[6][5] ),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05787_ (.A1(_00708_),
    .A2(_00795_),
    .B(_00797_),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05788_ (.I(_00798_),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05789_ (.I(net201),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05790_ (.I(\as2650.debug_psl[4] ),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05791_ (.I(\as2650.regs[0][5] ),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05792_ (.A1(_00715_),
    .A2(_00801_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05793_ (.A1(_00800_),
    .A2(\as2650.regs[4][5] ),
    .B(_00802_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05794_ (.I0(_00788_),
    .I1(_00794_),
    .I2(_00799_),
    .I3(_00803_),
    .S0(_00735_),
    .S1(_00768_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05795_ (.I(_00804_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05796_ (.A1(_00779_),
    .A2(_00617_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05797_ (.A1(_00743_),
    .A2(_00780_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05798_ (.A1(_00743_),
    .A2(\as2650.instruction_args_latch[5] ),
    .B1(_00806_),
    .B2(_00807_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05799_ (.A1(_00662_),
    .A2(_00805_),
    .B(_00808_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05800_ (.I(_00809_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05801_ (.I(_00657_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05802_ (.I(\as2650.regs[3][3] ),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05803_ (.A1(_00796_),
    .A2(\as2650.regs[7][3] ),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05804_ (.A1(_00708_),
    .A2(_00812_),
    .B(_00813_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05805_ (.I0(\as2650.regs[1][3] ),
    .I1(\as2650.regs[5][3] ),
    .S(_00800_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05806_ (.I(_00815_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05807_ (.I(_00816_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05808_ (.I(\as2650.regs[2][3] ),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05809_ (.A1(_00707_),
    .A2(\as2650.regs[6][3] ),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05810_ (.A1(_00796_),
    .A2(_00818_),
    .B(_00819_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05811_ (.I(_00820_),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05812_ (.I(\as2650.regs[0][3] ),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05813_ (.A1(_00753_),
    .A2(_00821_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05814_ (.A1(_00789_),
    .A2(\as2650.regs[4][3] ),
    .B(_00822_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05815_ (.I(_00823_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05816_ (.I(_00824_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05817_ (.I(_00825_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05818_ (.I(_00826_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05819_ (.I0(_00814_),
    .I1(_00817_),
    .I2(net198),
    .I3(_00827_),
    .S0(_00734_),
    .S1(_00704_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05820_ (.A1(_00811_),
    .A2(\as2650.instruction_args_latch[3] ),
    .A3(_00749_),
    .A4(_00828_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05821_ (.I(_00814_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _05822_ (.I(_00817_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05823_ (.I(net198),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05824_ (.I(_00823_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05825_ (.I0(_00830_),
    .I1(_00831_),
    .I2(_00832_),
    .I3(_00833_),
    .S0(_00734_),
    .S1(_00704_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05826_ (.A1(\as2650.indirect_target[3] ),
    .A2(_00621_),
    .B1(_00623_),
    .B2(\as2650.PC[3] ),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05827_ (.I(_00609_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05828_ (.A1(net305),
    .A2(_00836_),
    .A3(_00612_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05829_ (.A1(_00835_),
    .A2(_00837_),
    .B(_00657_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05830_ (.A1(_00811_),
    .A2(\as2650.instruction_args_latch[3] ),
    .B1(_00613_),
    .B2(_00838_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05831_ (.A1(_00661_),
    .A2(_00834_),
    .B(_00839_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05832_ (.A1(_00829_),
    .A2(_00840_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05833_ (.I(\as2650.regs[3][0] ),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05834_ (.A1(_00707_),
    .A2(\as2650.regs[7][0] ),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05835_ (.A1(_00692_),
    .A2(_00842_),
    .B(_00843_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05836_ (.I(_00789_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05837_ (.I0(\as2650.regs[1][0] ),
    .I1(\as2650.regs[5][0] ),
    .S(_00845_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05838_ (.I(_00723_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05839_ (.I(\as2650.regs[2][0] ),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05840_ (.A1(_00724_),
    .A2(\as2650.regs[6][0] ),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05841_ (.A1(_00847_),
    .A2(_00848_),
    .B(_00849_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05842_ (.I(_00850_),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05843_ (.I(\as2650.regs[0][0] ),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05844_ (.A1(_00753_),
    .A2(_00851_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05845_ (.A1(_00715_),
    .A2(\as2650.regs[4][0] ),
    .B(_00852_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05846_ (.I(_00853_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05847_ (.I(_00854_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05848_ (.I(_00855_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05849_ (.I0(_00844_),
    .I1(_00846_),
    .I2(net195),
    .I3(_00856_),
    .S0(net346),
    .S1(_00703_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05850_ (.A1(\as2650.instruction_args_latch[0] ),
    .A2(_00742_),
    .A3(_00659_),
    .A4(_00857_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05851_ (.A1(_00588_),
    .A2(_00658_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05852_ (.I(\as2650.regs[3][1] ),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05853_ (.A1(_00724_),
    .A2(\as2650.regs[7][1] ),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05854_ (.A1(_00847_),
    .A2(_00860_),
    .B(_00861_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05855_ (.I(\as2650.regs[5][1] ),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05856_ (.A1(_00723_),
    .A2(_00863_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05857_ (.A1(_00845_),
    .A2(\as2650.regs[1][1] ),
    .B(_00864_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05858_ (.I(_00865_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05859_ (.I(\as2650.regs[2][1] ),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05860_ (.A1(_00723_),
    .A2(\as2650.regs[6][1] ),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05861_ (.A1(_00845_),
    .A2(_00867_),
    .B(_00868_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05862_ (.I(_00869_),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05863_ (.I(\as2650.regs[0][1] ),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05864_ (.A1(_00689_),
    .A2(_00870_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05865_ (.A1(_00715_),
    .A2(\as2650.regs[4][1] ),
    .B(_00871_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05866_ (.I(_00872_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05867_ (.I(_00873_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05868_ (.I(_00874_),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05869_ (.I0(_00862_),
    .I1(_00866_),
    .I2(net196),
    .I3(_00875_),
    .S0(net345),
    .S1(_00702_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05870_ (.A1(net305),
    .A2(_00836_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05871_ (.A1(_00588_),
    .A2(\as2650.instruction_args_latch[1] ),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05872_ (.A1(_00657_),
    .A2(_00877_),
    .B(_00878_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05873_ (.A1(_00859_),
    .A2(_00876_),
    .B(_00879_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05874_ (.I(_00876_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05875_ (.A1(_00859_),
    .A2(_00881_),
    .A3(_00879_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05876_ (.A1(_00858_),
    .A2(_00880_),
    .B(_00882_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05877_ (.I(\as2650.regs[3][2] ),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05878_ (.A1(_00707_),
    .A2(\as2650.regs[7][2] ),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05879_ (.A1(_00692_),
    .A2(_00884_),
    .B(_00885_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05880_ (.I0(\as2650.regs[1][2] ),
    .I1(\as2650.regs[5][2] ),
    .S(_00800_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05881_ (.I(_00887_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05882_ (.I(_00888_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05883_ (.I(\as2650.regs[2][2] ),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05884_ (.A1(_00845_),
    .A2(\as2650.regs[6][2] ),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05885_ (.A1(_00847_),
    .A2(_00890_),
    .B(_00891_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05886_ (.I(_00892_),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05887_ (.I(\as2650.regs[0][2] ),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05888_ (.A1(_00689_),
    .A2(_00893_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05889_ (.A1(_00800_),
    .A2(\as2650.regs[4][2] ),
    .B(_00894_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05890_ (.I(_00895_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05891_ (.I(_00896_),
    .Z(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05892_ (.I(_00897_),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05893_ (.I0(_00886_),
    .I1(_00889_),
    .I2(net197),
    .I3(_00898_),
    .S0(net345),
    .S1(_00703_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _05894_ (.A1(_00742_),
    .A2(\as2650.instruction_args_latch[2] ),
    .A3(_00659_),
    .A4(_00899_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05895_ (.A1(net305),
    .A2(_00836_),
    .B(_00612_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05896_ (.A1(_00589_),
    .A2(_00837_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05897_ (.A1(_00901_),
    .A2(_00902_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _05898_ (.A1(_00742_),
    .A2(\as2650.instruction_args_latch[2] ),
    .B1(_00859_),
    .B2(_00899_),
    .C(_00903_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05899_ (.A1(_00904_),
    .A2(_00900_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05900_ (.A1(_00883_),
    .A2(_00905_),
    .B(_00900_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05901_ (.A1(_00841_),
    .A2(_00906_),
    .B(_00829_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05902_ (.I(\as2650.regs[3][4] ),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05903_ (.A1(_00796_),
    .A2(\as2650.regs[7][4] ),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05904_ (.A1(_00708_),
    .A2(_00908_),
    .B(_00909_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05905_ (.I(_00910_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05906_ (.I0(\as2650.regs[1][4] ),
    .I1(\as2650.regs[5][4] ),
    .S(_00789_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05907_ (.I(_00912_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05908_ (.I(_00913_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _05909_ (.I(_00914_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05910_ (.I(\as2650.regs[2][4] ),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05911_ (.A1(_00847_),
    .A2(\as2650.regs[6][4] ),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05912_ (.A1(_00692_),
    .A2(_00916_),
    .B(_00917_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05913_ (.I(_00918_),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05914_ (.I(net200),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05915_ (.I(\as2650.regs[0][4] ),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05916_ (.A1(_00753_),
    .A2(_00920_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05917_ (.A1(_00690_),
    .A2(\as2650.regs[4][4] ),
    .B(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05918_ (.I(_00922_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05919_ (.I0(_00911_),
    .I1(_00915_),
    .I2(_00919_),
    .I3(_00923_),
    .S0(_00734_),
    .S1(_00703_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05920_ (.A1(_00660_),
    .A2(_00924_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05921_ (.A1(_00613_),
    .A2(_00616_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05922_ (.A1(_00779_),
    .A2(_00926_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05923_ (.A1(_00811_),
    .A2(\as2650.instruction_args_latch[4] ),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05924_ (.A1(_00811_),
    .A2(_00927_),
    .B(_00928_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05925_ (.A1(_00925_),
    .A2(_00929_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05926_ (.A1(_00661_),
    .A2(_00804_),
    .A3(_00808_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05927_ (.A1(_00925_),
    .A2(_00929_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05928_ (.I(_00932_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05929_ (.A1(_00907_),
    .A2(_00930_),
    .B(_00931_),
    .C(_00933_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05930_ (.I0(_00697_),
    .I1(_00720_),
    .I2(net203),
    .I3(_00729_),
    .S0(_00735_),
    .S1(_00768_),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05931_ (.A1(_00744_),
    .A2(\as2650.instruction_args_latch[7] ),
    .A3(_00749_),
    .A4(_00935_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05932_ (.A1(_00770_),
    .A2(_00936_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05933_ (.A1(_00784_),
    .A2(_00810_),
    .A3(_00934_),
    .B(_00937_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05934_ (.I(_00938_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05935_ (.I(_00625_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05936_ (.A1(_00940_),
    .A2(_00627_),
    .B(_00629_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05937_ (.A1(_00744_),
    .A2(_00630_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05938_ (.A1(_00745_),
    .A2(\as2650.instruction_args_latch[11] ),
    .B1(_00941_),
    .B2(_00942_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05939_ (.I(_00748_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05940_ (.A1(_00740_),
    .A2(_00622_),
    .B(_00624_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05941_ (.A1(_00589_),
    .A2(_00940_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05942_ (.A1(_00944_),
    .A2(\as2650.instruction_args_latch[9] ),
    .B1(_00945_),
    .B2(_00946_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05943_ (.A1(_00740_),
    .A2(_00622_),
    .B(_00589_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05944_ (.A1(_00740_),
    .A2(_00622_),
    .B(_00948_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05945_ (.A1(_00944_),
    .A2(\as2650.instruction_args_latch[8] ),
    .B(_00949_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05946_ (.A1(_00940_),
    .A2(_00627_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05947_ (.A1(_00940_),
    .A2(_00627_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05948_ (.A1(_00944_),
    .A2(_00952_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05949_ (.A1(_00745_),
    .A2(\as2650.instruction_args_latch[10] ),
    .B1(_00951_),
    .B2(_00953_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05950_ (.A1(_00943_),
    .A2(_00947_),
    .A3(_00950_),
    .A4(_00954_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _05951_ (.A1(_00747_),
    .A2(_00939_),
    .A3(_00955_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05952_ (.A1(_00645_),
    .A2(\as2650.extend ),
    .B(\as2650.instruction_args_latch[13] ),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05953_ (.I(\as2650.page_reg[0] ),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05954_ (.A1(_00958_),
    .A2(_00646_),
    .B(_00590_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05955_ (.A1(_00633_),
    .A2(_00637_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05956_ (.A1(_00957_),
    .A2(_00959_),
    .B1(_00960_),
    .B2(_00590_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05957_ (.A1(_00630_),
    .A2(_00632_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05958_ (.A1(_00744_),
    .A2(\as2650.instruction_args_latch[12] ),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _05959_ (.A1(_00944_),
    .A2(_00633_),
    .A3(_00962_),
    .B(_00963_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05960_ (.A1(_00961_),
    .A2(_00964_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05961_ (.A1(_00656_),
    .A2(_00956_),
    .A3(_00965_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05962_ (.A1(_00651_),
    .A2(_00966_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05963_ (.I(_00967_),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05964_ (.A1(net227),
    .A2(net246),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05965_ (.I(_00968_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05966_ (.A1(_00747_),
    .A2(net429),
    .A3(_00955_),
    .A4(_00965_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05967_ (.A1(_00656_),
    .A2(_00970_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05968_ (.I(_00971_),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05969_ (.A1(net226),
    .A2(net245),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05970_ (.I(_00747_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05971_ (.I(_00950_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05972_ (.A1(_00947_),
    .A2(_00974_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05973_ (.I(_00954_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05974_ (.A1(_00973_),
    .A2(_00939_),
    .A3(_00975_),
    .A4(_00976_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05975_ (.A1(_00943_),
    .A2(_00977_),
    .B(_00956_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05976_ (.I(_00978_),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05977_ (.A1(net223),
    .A2(net242),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05978_ (.I(net236),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05979_ (.I(_00947_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05980_ (.I(_00973_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05981_ (.I(_00939_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05982_ (.I(_00974_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05983_ (.A1(_00982_),
    .A2(_00983_),
    .A3(_00984_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05984_ (.A1(_00982_),
    .A2(_00983_),
    .A3(_00975_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05985_ (.A1(_00981_),
    .A2(_00985_),
    .B(_00986_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05986_ (.I(_00987_),
    .ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05987_ (.A1(_00973_),
    .A2(_00939_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _05988_ (.A1(net235),
    .A2(_00988_),
    .A3(_00974_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _05989_ (.A1(net224),
    .A2(_00956_),
    .A3(_00964_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05990_ (.A1(_00980_),
    .A2(net255),
    .B(_00989_),
    .C(_00990_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05991_ (.A1(_00982_),
    .A2(_00983_),
    .A3(_00975_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _05992_ (.A1(net222),
    .A2(_00976_),
    .A3(_00992_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _05993_ (.A1(_00973_),
    .A2(_00983_),
    .A3(_00955_),
    .A4(_00964_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _05994_ (.A1(net225),
    .A2(_00961_),
    .A3(_00994_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05995_ (.A1(net236),
    .A2(_00987_),
    .B(_00993_),
    .C(_00995_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05996_ (.A1(_00972_),
    .A2(_00979_),
    .A3(_00991_),
    .A4(_00996_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05997_ (.I(_00997_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05998_ (.A1(_00969_),
    .A2(_00998_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05999_ (.A1(\as2650.cycle[2] ),
    .A2(\as2650.cycle[8] ),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06000_ (.I(_00591_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06001_ (.I(\as2650.is_interrupt_cycle ),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06002_ (.A1(_01001_),
    .A2(_01002_),
    .A3(_00603_),
    .A4(_00596_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06003_ (.A1(_01000_),
    .A2(_01003_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06004_ (.A1(_00999_),
    .A2(_01004_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06005_ (.I(_01005_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06006_ (.I(_01006_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06007_ (.I(_01007_),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06008_ (.A1(_00961_),
    .A2(_00994_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06009_ (.I(_01008_),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06010_ (.A1(_00956_),
    .A2(_00964_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06011_ (.I(_01009_),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06012_ (.A1(_00976_),
    .A2(_00992_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06013_ (.I(_01010_),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06014_ (.A1(_00988_),
    .A2(_00974_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06015_ (.I(_01011_),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06016_ (.I(_00721_),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06017_ (.I(_00758_),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06018_ (.I(_00793_),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06019_ (.I(_00914_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06020_ (.I(_01012_),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06021_ (.I(_00816_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06022_ (.I(_01013_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06023_ (.I(_01014_),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06024_ (.I(_00889_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06025_ (.I(_01015_),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06026_ (.I(_00866_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06027_ (.I(_01016_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06028_ (.I(_01017_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06029_ (.I(_01018_),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06030_ (.I(_00846_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06031_ (.I(_01019_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06032_ (.I(_01020_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06033_ (.I(_01021_),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06034_ (.I(_00730_),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06035_ (.I(_00767_),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06036_ (.I(_00803_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06037_ (.I(_01022_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06038_ (.I(_01023_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06039_ (.I(_01024_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06040_ (.I(_01025_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06041_ (.I(_01026_),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06042_ (.I(_00922_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06043_ (.I(_01027_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06044_ (.I(_01028_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06045_ (.I(_01029_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06046_ (.I(_01030_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06047_ (.I(_01031_),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06048_ (.A1(wb_reset_override),
    .A2(wb_reset_override_en),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06049_ (.A1(wb_reset_override_en),
    .A2(net33),
    .B(_01032_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06050_ (.A1(net66),
    .A2(_01033_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06051_ (.I(_01034_),
    .ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06052_ (.A1(_00982_),
    .A2(_00936_),
    .ZN(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06053_ (.A1(_00784_),
    .A2(_00810_),
    .A3(net348),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06054_ (.A1(_00770_),
    .A2(_01036_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06055_ (.A1(_01035_),
    .A2(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06056_ (.I(_01038_),
    .ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06057_ (.A1(net234),
    .A2(_01038_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06058_ (.I(\as2650.instruction_args_latch[0] ),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06059_ (.I(_00745_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06060_ (.A1(_01040_),
    .A2(_01041_),
    .A3(_00749_),
    .A4(_00857_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06061_ (.I(_00859_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06062_ (.I(_01043_),
    .Z(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06063_ (.A1(\as2650.PC[0] ),
    .A2(_00641_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06064_ (.A1(\as2650.indirect_target[0] ),
    .A2(_00635_),
    .B1(_00594_),
    .B2(\as2650.cycle[4] ),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06065_ (.A1(_01045_),
    .A2(_01046_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06066_ (.A1(_01041_),
    .A2(_00836_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06067_ (.A1(_01040_),
    .A2(_01041_),
    .B1(_01044_),
    .B2(_00857_),
    .C1(_01047_),
    .C2(_01048_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06068_ (.A1(_01042_),
    .A2(_01049_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06069_ (.A1(net221),
    .A2(_01050_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06070_ (.A1(_01043_),
    .A2(_00881_),
    .A3(_00879_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06071_ (.A1(_01052_),
    .A2(_00858_),
    .A3(_00880_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06072_ (.A1(_01052_),
    .A2(_00880_),
    .B(_00858_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06073_ (.A1(_01053_),
    .A2(_01054_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06074_ (.A1(net228),
    .A2(_01055_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06075_ (.A1(_00883_),
    .A2(_00905_),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06076_ (.I(_01057_),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06077_ (.A1(net229),
    .A2(net248),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06078_ (.A1(_00841_),
    .A2(net353),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06079_ (.I(_01059_),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06080_ (.I(net249),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06081_ (.A1(net230),
    .A2(_01060_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06082_ (.A1(_01051_),
    .A2(_01056_),
    .A3(_01058_),
    .A4(_01061_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06083_ (.A1(net350),
    .A2(_00930_),
    .Z(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06084_ (.I(_01063_),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06085_ (.A1(net231),
    .A2(net250),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06086_ (.A1(net349),
    .A2(_00930_),
    .B(_00933_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06087_ (.A1(_00810_),
    .A2(_00931_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06088_ (.A1(_01065_),
    .A2(_01066_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06089_ (.I(_01067_),
    .ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06090_ (.A1(net232),
    .A2(net251),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06091_ (.A1(_00810_),
    .A2(_00934_),
    .B(_00784_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06092_ (.A1(_01036_),
    .A2(_01069_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06093_ (.I(_01070_),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06094_ (.A1(net233),
    .A2(net252),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06095_ (.A1(_01062_),
    .A2(_01064_),
    .A3(_01068_),
    .A4(_01071_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06096_ (.A1(net234),
    .A2(_01038_),
    .Z(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06097_ (.A1(_01039_),
    .A2(_01072_),
    .A3(_01073_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06098_ (.I(_01074_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06099_ (.A1(_00999_),
    .A2(_01000_),
    .A3(_01003_),
    .A4(_01075_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06100_ (.I(_01076_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06101_ (.I(_01077_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06102_ (.I(_01078_),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06103_ (.I(_01055_),
    .ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06104_ (.I(_01050_),
    .ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06105_ (.I(_00666_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06106_ (.I(_01079_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06107_ (.I(_01080_),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _06108_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(net256),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06109_ (.I(_01081_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06110_ (.I(_01082_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06111_ (.I(_01083_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06112_ (.I(_01084_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06113_ (.I(_01085_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06114_ (.I(_01086_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06115_ (.I(_01087_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06116_ (.I(\as2650.cycle[11] ),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06117_ (.A1(net48),
    .A2(net47),
    .A3(net49),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06118_ (.A1(net44),
    .A2(net43),
    .A3(net46),
    .A4(net45),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06119_ (.I(\as2650.debug_psu[5] ),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06120_ (.A1(_01090_),
    .A2(_01091_),
    .B(_01092_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06121_ (.I(_01093_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06122_ (.I(_00700_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06123_ (.I(_01095_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06124_ (.I(_01096_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06125_ (.I(_01097_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06126_ (.A1(_01098_),
    .A2(_00969_),
    .A3(_00998_),
    .A4(_01075_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06127_ (.I(_01099_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06128_ (.I(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06129_ (.I(_01101_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06130_ (.I(\as2650.extend ),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06131_ (.I(_00669_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06132_ (.I(_00671_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06133_ (.I(_00673_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06134_ (.I(net40),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06135_ (.A1(_01104_),
    .A2(_01105_),
    .A3(_01106_),
    .B(_01107_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _06136_ (.A1(_01104_),
    .A2(net52),
    .A3(_00671_),
    .A4(_00673_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06137_ (.A1(_01108_),
    .A2(_01109_),
    .B(_00666_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06138_ (.I(_00665_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06139_ (.A1(net60),
    .A2(_01111_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06140_ (.A1(\as2650.insin[2] ),
    .A2(_00700_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06141_ (.A1(_00700_),
    .A2(_01110_),
    .A3(_01112_),
    .B(_01113_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06142_ (.I(_01114_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06143_ (.A1(_01103_),
    .A2(_01115_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06144_ (.I(_00664_),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _06145_ (.A1(_01104_),
    .A2(net53),
    .A3(_01105_),
    .A4(_01106_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06146_ (.I(_01104_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06147_ (.I(net41),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06148_ (.A1(_01119_),
    .A2(_01105_),
    .A3(_01106_),
    .B(_01120_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06149_ (.A1(_01118_),
    .A2(_01121_),
    .B(_01079_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06150_ (.A1(net61),
    .A2(_01111_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06151_ (.A1(_01122_),
    .A2(_01123_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06152_ (.A1(_01117_),
    .A2(_01124_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06153_ (.A1(\as2650.insin[3] ),
    .A2(_01095_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06154_ (.A1(_01125_),
    .A2(_01126_),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06155_ (.A1(_01116_),
    .A2(_01127_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06156_ (.I(_01103_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06157_ (.I(_01129_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06158_ (.I(_01130_),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06159_ (.A1(_01119_),
    .A2(_01105_),
    .A3(_01106_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06160_ (.I(_01132_),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06161_ (.I(net57),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06162_ (.A1(_01134_),
    .A2(_01133_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06163_ (.A1(net36),
    .A2(_01133_),
    .B(_01135_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06164_ (.A1(net65),
    .A2(_01080_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06165_ (.A1(_01080_),
    .A2(_01136_),
    .B(_01137_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06166_ (.A1(_00664_),
    .A2(_01138_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06167_ (.A1(\as2650.insin[7] ),
    .A2(_01096_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06168_ (.A1(_01139_),
    .A2(_01140_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06169_ (.I(_01141_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06170_ (.I(net56),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06171_ (.A1(_01143_),
    .A2(_01132_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06172_ (.A1(net35),
    .A2(_01133_),
    .B(_01144_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06173_ (.A1(net64),
    .A2(_01079_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06174_ (.A1(_01079_),
    .A2(_01145_),
    .B(_01146_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06175_ (.A1(_00664_),
    .A2(_01147_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06176_ (.A1(\as2650.insin[6] ),
    .A2(_01095_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06177_ (.A1(_01148_),
    .A2(_01149_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06178_ (.I(_01150_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06179_ (.A1(_01142_),
    .A2(_01151_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06180_ (.I(_01111_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06181_ (.I(_01132_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06182_ (.I(net55),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06183_ (.A1(_01155_),
    .A2(_01154_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06184_ (.A1(net34),
    .A2(_01154_),
    .B(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06185_ (.A1(_01111_),
    .A2(_01157_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06186_ (.A1(net63),
    .A2(_01153_),
    .B(_01158_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06187_ (.I(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06188_ (.A1(\as2650.insin[5] ),
    .A2(_01097_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06189_ (.A1(_01097_),
    .A2(_01160_),
    .B(_01161_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06190_ (.I(_01162_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06191_ (.A1(_01148_),
    .A2(_01149_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06192_ (.I(_01164_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06193_ (.A1(_01142_),
    .A2(_01165_),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06194_ (.I(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06195_ (.A1(_01163_),
    .A2(_01167_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06196_ (.I(_01168_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06197_ (.I(_01115_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06198_ (.I(_01127_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06199_ (.A1(_01170_),
    .A2(_01171_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06200_ (.A1(\as2650.insin[4] ),
    .A2(_01096_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06201_ (.I(net54),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06202_ (.A1(_01174_),
    .A2(_01133_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06203_ (.A1(net42),
    .A2(_01154_),
    .B(_01175_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06204_ (.A1(net62),
    .A2(_01080_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06205_ (.A1(net139),
    .A2(_01176_),
    .B(_01177_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06206_ (.A1(_01117_),
    .A2(_01178_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06207_ (.A1(_01173_),
    .A2(_01179_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06208_ (.I(_01180_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06209_ (.A1(_01130_),
    .A2(_01172_),
    .A3(_01181_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06210_ (.I(_01182_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06211_ (.A1(_01152_),
    .A2(_01169_),
    .B(_01183_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06212_ (.I(_00736_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06213_ (.I(_01185_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06214_ (.I(_00706_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06215_ (.I(_01187_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06216_ (.A1(_01186_),
    .A2(_01188_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06217_ (.I(_01172_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06218_ (.I(_01190_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06219_ (.A1(_01103_),
    .A2(_01180_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06220_ (.I(_01192_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06221_ (.A1(_01191_),
    .A2(_01193_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06222_ (.I(_01162_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06223_ (.A1(_01139_),
    .A2(_01140_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06224_ (.A1(_01196_),
    .A2(_01151_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06225_ (.I(_01197_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06226_ (.A1(_01195_),
    .A2(_01198_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06227_ (.I(_01199_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06228_ (.A1(_01194_),
    .A2(_01200_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06229_ (.A1(_01189_),
    .A2(_01201_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06230_ (.I(_01103_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06231_ (.I(_01203_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06232_ (.A1(_01173_),
    .A2(_01179_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06233_ (.A1(_01205_),
    .A2(_01195_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06234_ (.A1(_01196_),
    .A2(_01164_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06235_ (.A1(_01204_),
    .A2(_01191_),
    .A3(_01206_),
    .A4(_01207_),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06236_ (.A1(_01095_),
    .A2(_01122_),
    .A3(_01123_),
    .B(_01126_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06237_ (.A1(_01115_),
    .A2(_01209_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06238_ (.I(_01210_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06239_ (.I(_01211_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06240_ (.I(_01212_),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06241_ (.I(_01213_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06242_ (.I(_01214_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06243_ (.I(_01215_),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06244_ (.A1(_01115_),
    .A2(_01209_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06245_ (.A1(_01208_),
    .A2(_01216_),
    .A3(_01217_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06246_ (.A1(_01184_),
    .A2(_01202_),
    .A3(_01218_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06247_ (.A1(_01131_),
    .A2(_01219_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06248_ (.A1(_01128_),
    .A2(_01220_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06249_ (.I(_01221_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06250_ (.A1(_01102_),
    .A2(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06251_ (.I(_00688_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06252_ (.I(_01210_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06253_ (.I(_01225_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06254_ (.I(_01226_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06255_ (.A1(_01186_),
    .A2(_01227_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06256_ (.A1(_01129_),
    .A2(_01224_),
    .A3(_01228_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06257_ (.A1(_01142_),
    .A2(_01165_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06258_ (.I(_01230_),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06259_ (.A1(_01206_),
    .A2(_01229_),
    .A3(_01231_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06260_ (.I(_01232_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06261_ (.A1(_01089_),
    .A2(_01223_),
    .A3(_01233_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06262_ (.A1(_01089_),
    .A2(_01094_),
    .B(_01234_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06263_ (.A1(_01088_),
    .A2(_01235_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06264_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(net355),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06265_ (.I(_01236_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06266_ (.I(_01237_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06267_ (.I(_01238_),
    .Z(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06268_ (.I(_01239_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06269_ (.I(_01240_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06270_ (.A1(_00969_),
    .A2(_00998_),
    .A3(_01075_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06271_ (.I(_01242_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06272_ (.I(_01243_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06273_ (.A1(_01098_),
    .A2(_01244_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06274_ (.A1(\as2650.cycle[11] ),
    .A2(_01245_),
    .B(_01093_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06275_ (.I(_01246_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06276_ (.A1(_01241_),
    .A2(_01247_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06277_ (.I(\as2650.cycle[4] ),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06278_ (.I(_01249_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06279_ (.I(_01250_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06280_ (.I(_01251_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06281_ (.A1(_00999_),
    .A2(_01039_),
    .A3(net351),
    .A4(_01073_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06282_ (.I(_01253_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06283_ (.I(_01254_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06284_ (.I(_01255_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06285_ (.I(_01253_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06286_ (.I(_01257_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06287_ (.I(_01258_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06288_ (.A1(_00645_),
    .A2(_01128_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06289_ (.I(_01260_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06290_ (.I(\as2650.cycle[6] ),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06291_ (.I(_01262_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06292_ (.I(_01263_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06293_ (.I(_01264_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06294_ (.I(\as2650.relative_cyc ),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06295_ (.A1(_01266_),
    .A2(_01190_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06296_ (.I(_01267_),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06297_ (.A1(_01265_),
    .A2(_01268_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06298_ (.A1(_01259_),
    .A2(_01261_),
    .A3(_01269_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06299_ (.A1(_01252_),
    .A2(_01256_),
    .B(_01270_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06300_ (.A1(_01248_),
    .A2(_01271_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06301_ (.A1(_01192_),
    .A2(_01163_),
    .A3(_01213_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06302_ (.I(_01272_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06303_ (.I(_01100_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06304_ (.I(_01274_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06305_ (.I(_00680_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06306_ (.I(_01205_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06307_ (.I(_01277_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06308_ (.A1(_01096_),
    .A2(_01159_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06309_ (.A1(\as2650.insin[5] ),
    .A2(_01097_),
    .B(_01279_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06310_ (.I(_01280_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06311_ (.I(_01281_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06312_ (.I(_01282_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06313_ (.A1(_01278_),
    .A2(_01283_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06314_ (.A1(_01167_),
    .A2(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06315_ (.A1(_01131_),
    .A2(_01276_),
    .A3(_01216_),
    .A4(_01285_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06316_ (.I(_01286_),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06317_ (.A1(_01275_),
    .A2(_01287_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06318_ (.A1(_01248_),
    .A2(_01273_),
    .A3(_01288_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06319_ (.A1(_01240_),
    .A2(_01246_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06320_ (.I(_01289_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06321_ (.A1(\as2650.cycle[5] ),
    .A2(_01290_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06322_ (.I(_01291_),
    .Z(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06323_ (.I(_01041_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06324_ (.I(_01292_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06325_ (.I(_01244_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06326_ (.I(_01294_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06327_ (.A1(_01171_),
    .A2(_01181_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06328_ (.I(_01296_),
    .Z(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06329_ (.I(_01297_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06330_ (.I(\as2650.instruction_args_latch[15] ),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06331_ (.I(_01209_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06332_ (.A1(_00647_),
    .A2(_01300_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06333_ (.A1(_01299_),
    .A2(_01301_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06334_ (.A1(_01249_),
    .A2(_01302_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06335_ (.I(_01243_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06336_ (.I(_01304_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06337_ (.I(_01305_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06338_ (.I(_01098_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06339_ (.A1(_01307_),
    .A2(_01287_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06340_ (.A1(_01298_),
    .A2(_01303_),
    .B(_01306_),
    .C(_01308_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06341_ (.A1(_01293_),
    .A2(_01295_),
    .B(_01289_),
    .C(_01309_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06342_ (.I(_01310_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06343_ (.A1(\as2650.cycle[7] ),
    .A2(_01290_),
    .Z(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06344_ (.I(_01311_),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06345_ (.A1(\as2650.cycle[2] ),
    .A2(_01290_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06346_ (.I(_01312_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06347_ (.I(\as2650.cycle[1] ),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06348_ (.A1(_01313_),
    .A2(_01248_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06349_ (.I(\as2650.cycle[6] ),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06350_ (.I(_01314_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06351_ (.I(_01268_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06352_ (.A1(_01138_),
    .A2(_01301_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06353_ (.A1(_01170_),
    .A2(_01317_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06354_ (.I(_01318_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06355_ (.I(_01319_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06356_ (.A1(\as2650.cycle[11] ),
    .A2(_01245_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06357_ (.A1(_01170_),
    .A2(_01171_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06358_ (.A1(_01317_),
    .A2(_01322_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06359_ (.I(_01323_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06360_ (.A1(_01181_),
    .A2(_01324_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06361_ (.I(_01325_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06362_ (.A1(_01321_),
    .A2(_01322_),
    .B(_01326_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06363_ (.A1(_01261_),
    .A2(_01327_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06364_ (.A1(_01320_),
    .A2(_01328_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06365_ (.I(_01254_),
    .Z(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06366_ (.A1(_01316_),
    .A2(_01329_),
    .B(_01330_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06367_ (.I(_01250_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06368_ (.A1(_01299_),
    .A2(_01301_),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06369_ (.A1(_01332_),
    .A2(_01333_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06370_ (.I(_01334_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06371_ (.I(_01117_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06372_ (.I(_01287_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06373_ (.A1(_01205_),
    .A2(_01207_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06374_ (.I(_01338_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06375_ (.I(_01339_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06376_ (.A1(_01281_),
    .A2(_01339_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06377_ (.I(_01341_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06378_ (.I(_00935_),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06379_ (.I(_00778_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _06380_ (.I0(_00787_),
    .I1(net192),
    .I2(net201),
    .I3(_01025_),
    .S0(_01186_),
    .S1(_01188_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06381_ (.I(_01345_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06382_ (.I(_00924_),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06383_ (.I(_00834_),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06384_ (.I(_00899_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06385_ (.I(_00862_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06386_ (.I(_00865_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06387_ (.I(net196),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _06388_ (.I0(_01350_),
    .I1(_01351_),
    .I2(_01352_),
    .I3(_00872_),
    .S0(_00736_),
    .S1(_00706_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06389_ (.I(_00844_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06390_ (.I(_01021_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06391_ (.I(net195),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _06392_ (.I0(_01354_),
    .I1(_01355_),
    .I2(_01356_),
    .I3(_00853_),
    .S0(_01185_),
    .S1(_01187_),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06393_ (.A1(_01353_),
    .A2(_01357_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06394_ (.A1(_01349_),
    .A2(_01358_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06395_ (.A1(_01347_),
    .A2(_01348_),
    .A3(_01359_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06396_ (.A1(_01346_),
    .A2(_01360_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06397_ (.A1(_01344_),
    .A2(_01361_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06398_ (.A1(_01343_),
    .A2(_01362_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06399_ (.A1(_01141_),
    .A2(_01150_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06400_ (.A1(_01180_),
    .A2(_01364_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06401_ (.A1(_01280_),
    .A2(_01365_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06402_ (.I(_01366_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06403_ (.I(_00886_),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06404_ (.I(net206),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06405_ (.I(net189),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06406_ (.I(net197),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _06407_ (.I0(_01368_),
    .I1(_01369_),
    .I2(_01370_),
    .I3(_00895_),
    .S0(_01185_),
    .S1(_01187_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06408_ (.I(_00881_),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06409_ (.I(_00857_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06410_ (.A1(_01372_),
    .A2(_01373_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06411_ (.A1(_01371_),
    .A2(_01374_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06412_ (.A1(_00828_),
    .A2(_01375_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06413_ (.A1(_01347_),
    .A2(_01376_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06414_ (.A1(_01346_),
    .A2(_01377_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06415_ (.A1(_01344_),
    .A2(_01378_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06416_ (.A1(_01343_),
    .A2(_01379_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06417_ (.A1(_01367_),
    .A2(_01380_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06418_ (.A1(_00738_),
    .A2(_01340_),
    .B1(_01342_),
    .B2(_01363_),
    .C(_01381_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06419_ (.I(_01345_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06420_ (.A1(_01383_),
    .A2(_01360_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06421_ (.A1(_01346_),
    .A2(_01377_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06422_ (.A1(_01367_),
    .A2(_01385_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06423_ (.A1(_00805_),
    .A2(_01340_),
    .B1(_01341_),
    .B2(_01384_),
    .C(_01386_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06424_ (.I(_01347_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06425_ (.I(_00910_),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _06426_ (.I0(net208),
    .I1(net191),
    .I2(net200),
    .I3(_01031_),
    .S0(_01185_),
    .S1(_01187_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06427_ (.I(_01348_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06428_ (.A1(_01390_),
    .A2(_01359_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06429_ (.A1(_01389_),
    .A2(_01391_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06430_ (.A1(_01360_),
    .A2(_01392_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06431_ (.I(_01393_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06432_ (.A1(_01347_),
    .A2(_01376_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06433_ (.A1(_01367_),
    .A2(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06434_ (.A1(_01388_),
    .A2(_01340_),
    .B1(_01342_),
    .B2(_01394_),
    .C(_01396_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06435_ (.A1(_01162_),
    .A2(_01338_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06436_ (.A1(_01348_),
    .A2(_01375_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06437_ (.A1(_01162_),
    .A2(_01365_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06438_ (.I(_00828_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06439_ (.A1(_01401_),
    .A2(_01359_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06440_ (.A1(_01400_),
    .A2(_01402_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06441_ (.A1(_01390_),
    .A2(_01339_),
    .B1(_01398_),
    .B2(_01399_),
    .C(_01403_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06442_ (.I(_01371_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06443_ (.A1(_01405_),
    .A2(_01358_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06444_ (.A1(_01400_),
    .A2(_01406_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06445_ (.A1(_01405_),
    .A2(_01374_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06446_ (.A1(_01366_),
    .A2(_01408_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06447_ (.A1(_01405_),
    .A2(_01339_),
    .B(_01407_),
    .C(_01409_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06448_ (.I(_01373_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06449_ (.A1(_01411_),
    .A2(_01365_),
    .Z(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06450_ (.A1(_01358_),
    .A2(_01374_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06451_ (.A1(_01411_),
    .A2(_01365_),
    .B(_01366_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06452_ (.A1(_01413_),
    .A2(_01414_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06453_ (.A1(_01404_),
    .A2(_01410_),
    .A3(_01412_),
    .A4(_01415_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06454_ (.A1(_01387_),
    .A2(_01397_),
    .A3(_01416_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06455_ (.I(_01344_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06456_ (.I(_00769_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06457_ (.A1(_01419_),
    .A2(_01378_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06458_ (.A1(_01344_),
    .A2(_01361_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06459_ (.A1(_01342_),
    .A2(_01421_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06460_ (.A1(_01418_),
    .A2(_01340_),
    .B1(_01398_),
    .B2(_01420_),
    .C(_01422_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06461_ (.I(_01277_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06462_ (.A1(_01424_),
    .A2(_01165_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06463_ (.A1(_01382_),
    .A2(_01417_),
    .A3(_01423_),
    .B(_01425_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06464_ (.A1(_00680_),
    .A2(_01224_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06465_ (.A1(\as2650.debug_psl[6] ),
    .A2(_01188_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06466_ (.I(_01186_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06467_ (.A1(\as2650.debug_psl[7] ),
    .A2(_01429_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06468_ (.A1(_01428_),
    .A2(_01430_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06469_ (.A1(_01427_),
    .A2(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06470_ (.A1(_01278_),
    .A2(_01152_),
    .A3(_01432_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06471_ (.I(_01198_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06472_ (.A1(_01192_),
    .A2(_01434_),
    .A3(_01189_),
    .A4(_01322_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06473_ (.A1(_01192_),
    .A2(_01197_),
    .A3(_01189_),
    .A4(_01217_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06474_ (.I(_01436_),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06475_ (.I(_01437_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06476_ (.I(_01438_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06477_ (.A1(_01300_),
    .A2(_01424_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06478_ (.A1(_01434_),
    .A2(_01431_),
    .B(_01439_),
    .C(_01440_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _06479_ (.A1(_01426_),
    .A2(_01433_),
    .A3(_01435_),
    .A4(_01441_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06480_ (.I(_01442_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06481_ (.I(_01443_),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06482_ (.I(_01444_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06483_ (.A1(_01222_),
    .A2(_01445_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06484_ (.A1(_01336_),
    .A2(_01337_),
    .A3(_01446_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06485_ (.A1(_01335_),
    .A2(_01447_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06486_ (.I(_01254_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06487_ (.I(_01002_),
    .Z(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06488_ (.A1(_01315_),
    .A2(_01331_),
    .B1(_01448_),
    .B2(_01449_),
    .C(_01450_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06489_ (.A1(_01314_),
    .A2(_01253_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06490_ (.I(_01452_),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06491_ (.I(_01453_),
    .Z(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06492_ (.A1(_01260_),
    .A2(_01268_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06493_ (.I(_01455_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06494_ (.A1(_01089_),
    .A2(_01322_),
    .A3(_01456_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06495_ (.A1(_01247_),
    .A2(_01451_),
    .B1(_01454_),
    .B2(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06496_ (.A1(_01088_),
    .A2(_01458_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06497_ (.A1(_01266_),
    .A2(_01191_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06498_ (.A1(_01262_),
    .A2(_01459_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06499_ (.I(_01151_),
    .Z(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06500_ (.I(_01283_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06501_ (.A1(_01183_),
    .A2(_01461_),
    .A3(_01462_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06502_ (.A1(_01257_),
    .A2(_01460_),
    .A3(_01463_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06503_ (.I(_01464_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06504_ (.I(_01465_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06505_ (.A1(_01290_),
    .A2(_01466_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06506_ (.I(_01467_),
    .Z(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06507_ (.A1(_01264_),
    .A2(_01304_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06508_ (.I(_01468_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06509_ (.A1(_01089_),
    .A2(_01316_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06510_ (.A1(_01260_),
    .A2(_01267_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06511_ (.I(_01471_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06512_ (.A1(_01278_),
    .A2(_01323_),
    .A3(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06513_ (.I(_01473_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06514_ (.I(_01474_),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06515_ (.A1(_01463_),
    .A2(_01470_),
    .B1(_01475_),
    .B2(_01247_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06516_ (.I(\as2650.cycle[10] ),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06517_ (.A1(_01314_),
    .A2(_01267_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06518_ (.A1(\as2650.cycle[11] ),
    .A2(_01245_),
    .B(_01478_),
    .C(_01463_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06519_ (.I(_01117_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06520_ (.A1(_01233_),
    .A2(_01273_),
    .A3(_01287_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06521_ (.A1(_01446_),
    .A2(_01481_),
    .B(_01294_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06522_ (.A1(_01440_),
    .A2(_01303_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06523_ (.A1(_01480_),
    .A2(_01482_),
    .B(_01483_),
    .C(_01293_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06524_ (.A1(_01480_),
    .A2(_01305_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06525_ (.A1(_01479_),
    .A2(_01484_),
    .B(_01485_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06526_ (.A1(_01477_),
    .A2(\as2650.cycle[8] ),
    .A3(_01486_),
    .B(_01247_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06527_ (.I(_01241_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06528_ (.A1(_01469_),
    .A2(_01476_),
    .B(_01487_),
    .C(_01488_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06529_ (.I(_00856_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06530_ (.I(_01489_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06531_ (.I(_01490_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06532_ (.I(_01491_),
    .Z(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06533_ (.I(_01492_),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06534_ (.I(_00874_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06535_ (.I(_01493_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06536_ (.I(_01494_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06537_ (.I(_01495_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06538_ (.I(_01496_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06539_ (.I(_01497_),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06540_ (.I(_00897_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06541_ (.I(_01498_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06542_ (.I(_01499_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06543_ (.I(_01500_),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06544_ (.I(_00827_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06545_ (.I(_01501_),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06546_ (.I(wb_io3_test),
    .ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06547_ (.A1(_00969_),
    .A2(_00998_),
    .A3(_01075_),
    .A4(_01081_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06548_ (.I(_01502_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06549_ (.I(_01503_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06550_ (.I(_01504_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06551_ (.I(_01263_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06552_ (.A1(_01266_),
    .A2(_01506_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06553_ (.A1(_01203_),
    .A2(_01300_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06554_ (.A1(_00688_),
    .A2(_01228_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06555_ (.A1(_01203_),
    .A2(_01509_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06556_ (.A1(_01206_),
    .A2(_01207_),
    .A3(_01510_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06557_ (.A1(_01508_),
    .A2(_01511_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06558_ (.I(_01512_),
    .Z(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06559_ (.A1(_01001_),
    .A2(_01507_),
    .B(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06560_ (.A1(_01154_),
    .A2(_01505_),
    .A3(_01514_),
    .ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06561_ (.I(_01084_),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06562_ (.A1(_01515_),
    .A2(_01246_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06563_ (.I(_01516_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06564_ (.I(\as2650.io_bus_we ),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06565_ (.I(\as2650.ext_io_addr[7] ),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06566_ (.I(_01518_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06567_ (.I(\as2650.ext_io_addr[6] ),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06568_ (.I(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06569_ (.A1(_01517_),
    .A2(_01519_),
    .A3(_01521_),
    .ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06570_ (.I(_01519_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06571_ (.A1(\as2650.io_bus_we ),
    .A2(_01522_),
    .A3(_01521_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06572_ (.I(_01523_),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06573_ (.A1(_01517_),
    .A2(_01522_),
    .A3(_01521_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06574_ (.A1(\as2650.io_bus_we ),
    .A2(_01519_),
    .A3(_01521_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06575_ (.I(_01524_),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06576_ (.I(_01515_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06577_ (.I(_01525_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06578_ (.I(_01077_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06579_ (.I(_01196_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06580_ (.I(_01528_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06581_ (.A1(_01000_),
    .A2(_01529_),
    .A3(_01273_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06582_ (.I(_01530_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06583_ (.A1(_01529_),
    .A2(_01273_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06584_ (.A1(\as2650.cycle[2] ),
    .A2(_01532_),
    .B(_01514_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06585_ (.I(_01085_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06586_ (.A1(_01000_),
    .A2(_01255_),
    .B(_01533_),
    .C(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06587_ (.A1(net237),
    .A2(_01527_),
    .A3(_01531_),
    .A4(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06588_ (.A1(_01526_),
    .A2(_01536_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06589_ (.I(_01537_),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06590_ (.I(_01086_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06591_ (.A1(_01142_),
    .A2(_01272_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _06592_ (.A1(\as2650.cycle[2] ),
    .A2(\as2650.cycle[8] ),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06593_ (.A1(_01003_),
    .A2(_01306_),
    .B1(_01539_),
    .B2(_01540_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _06594_ (.A1(_01538_),
    .A2(_01514_),
    .A3(_01541_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06595_ (.I(_01542_),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06596_ (.I(_01005_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06597_ (.I(_01543_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06598_ (.I(_01544_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06599_ (.I(_01239_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06600_ (.I(_01546_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06601_ (.I(_01547_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06602_ (.A1(clknet_leaf_36_wb_clk_i),
    .A2(_01548_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06603_ (.A1(_01545_),
    .A2(clknet_1_0__leaf__01549_),
    .ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06604_ (.I(_01076_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06605_ (.I(_01550_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06606_ (.I(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06607_ (.A1(_01552_),
    .A2(clknet_1_1__leaf__01549_),
    .ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06608_ (.I(\web_behavior[0] ),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06609_ (.A1(\web_behavior[1] ),
    .A2(_01553_),
    .A3(clknet_leaf_149_wb_clk_i),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06610_ (.A1(\web_behavior[1] ),
    .A2(_01553_),
    .A3(clknet_leaf_149_wb_clk_i),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06611_ (.A1(net304),
    .A2(_01554_),
    .A3(_01555_),
    .ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06612_ (.I(wb_debug_carry),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06613_ (.I(\as2650.debug_psl[0] ),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06614_ (.I(_01557_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06615_ (.I(\as2650.debug_psl[6] ),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06616_ (.I(_01559_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06617_ (.I(wb_debug_cc),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06618_ (.A1(\as2650.insin[6] ),
    .A2(_01561_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06619_ (.A1(wb_debug_cc),
    .A2(_01560_),
    .B1(_01540_),
    .B2(_01562_),
    .C(_01556_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06620_ (.A1(_01556_),
    .A2(_01558_),
    .B(_01563_),
    .ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06621_ (.I(\as2650.debug_psl[7] ),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06622_ (.I(_01564_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06623_ (.A1(\as2650.insin[6] ),
    .A2(wb_debug_cc),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06624_ (.A1(wb_debug_cc),
    .A2(_01565_),
    .B1(_01540_),
    .B2(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06625_ (.I(\as2650.debug_psl[5] ),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06626_ (.I(_01568_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06627_ (.I(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06628_ (.A1(_01556_),
    .A2(_01570_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06629_ (.A1(_01556_),
    .A2(_01567_),
    .B(_01571_),
    .ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06630_ (.I(_00844_),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06631_ (.I(_00862_),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06632_ (.I(_00814_),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06633_ (.I(_00787_),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06634_ (.I(_00697_),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _06635_ (.A1(_01098_),
    .A2(_00968_),
    .A3(_00997_),
    .A4(_01074_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06636_ (.I(_01572_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06637_ (.I(_01573_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06638_ (.A1(_01277_),
    .A2(_01152_),
    .A3(_01282_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06639_ (.I(_01575_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06640_ (.I(_01224_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06641_ (.A1(_01129_),
    .A2(_01276_),
    .A3(_01577_),
    .A4(_01214_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06642_ (.A1(_01576_),
    .A2(_01578_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06643_ (.A1(_01574_),
    .A2(_01579_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06644_ (.A1(\as2650.chirp_ptr[1] ),
    .A2(\as2650.chirp_ptr[0] ),
    .A3(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06645_ (.A1(\as2650.chirp_ptr[2] ),
    .A2(_01581_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06646_ (.I(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06647_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01580_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06648_ (.A1(_01239_),
    .A2(_01584_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06649_ (.I(_01585_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06650_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01580_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06651_ (.A1(\as2650.chirp_ptr[1] ),
    .A2(_01586_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06652_ (.A1(_01239_),
    .A2(_01587_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06653_ (.I(_01588_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06654_ (.A1(_00178_),
    .A2(_00179_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06655_ (.A1(_01584_),
    .A2(_00179_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06656_ (.A1(_01589_),
    .A2(_01590_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06657_ (.A1(_01515_),
    .A2(_01583_),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06658_ (.I(_01592_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06659_ (.A1(_01583_),
    .A2(_00178_),
    .B1(_01591_),
    .B2(_00180_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06660_ (.I(_01592_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06661_ (.I(_01589_),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06662_ (.A1(_01593_),
    .A2(_01594_),
    .B(_01590_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06663_ (.A1(_01593_),
    .A2(_01587_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06664_ (.A1(_01593_),
    .A2(_01591_),
    .B(_01595_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06665_ (.I0(_01590_),
    .I1(_01594_),
    .S(_01592_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06666_ (.I(_01596_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06667_ (.A1(_01593_),
    .A2(_01594_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06668_ (.A1(_00180_),
    .A2(_01587_),
    .B(_01597_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06669_ (.I(_01357_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06670_ (.I(_01598_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06671_ (.I(_01531_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06672_ (.I(_01600_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06673_ (.I(_01006_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06674_ (.A1(net254),
    .A2(_01602_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06675_ (.I(_01543_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06676_ (.I(_01043_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06677_ (.I(_01605_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06678_ (.A1(_01043_),
    .A2(_01490_),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06679_ (.A1(_01606_),
    .A2(_01598_),
    .B(_01607_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06680_ (.A1(_01604_),
    .A2(_01608_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06681_ (.A1(_01603_),
    .A2(_01609_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06682_ (.A1(_01050_),
    .A2(_01551_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06683_ (.I(_01530_),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06684_ (.A1(_01551_),
    .A2(_01610_),
    .B(_01611_),
    .C(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06685_ (.A1(_01599_),
    .A2(_01601_),
    .B(_01613_),
    .ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06686_ (.I(_01353_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06687_ (.I(_01614_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06688_ (.I(_01615_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06689_ (.I(_01078_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06690_ (.A1(net255),
    .A2(_01007_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06691_ (.A1(_01044_),
    .A2(_01496_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06692_ (.A1(_01044_),
    .A2(_01353_),
    .B(_01619_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06693_ (.I(_01620_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06694_ (.A1(_01544_),
    .A2(_01621_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06695_ (.A1(_01618_),
    .A2(_01622_),
    .B(_01527_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06696_ (.A1(net247),
    .A2(_01617_),
    .B(_01612_),
    .C(_01623_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06697_ (.A1(_01616_),
    .A2(_01601_),
    .B(_01624_),
    .ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06698_ (.I(_01405_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06699_ (.I(_01625_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06700_ (.I(_01612_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06701_ (.I(_01550_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06702_ (.A1(net241),
    .A2(_01602_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06703_ (.A1(_01605_),
    .A2(net210),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06704_ (.A1(_01605_),
    .A2(_01371_),
    .B(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06705_ (.I(_01631_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06706_ (.A1(_01604_),
    .A2(_01632_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06707_ (.A1(_01629_),
    .A2(_01633_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06708_ (.A1(_01628_),
    .A2(_01634_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06709_ (.A1(net248),
    .A2(net238),
    .B(_01600_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06710_ (.A1(_01626_),
    .A2(_01627_),
    .B1(_01635_),
    .B2(_01636_),
    .ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06711_ (.I(_01390_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06712_ (.I(_01550_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06713_ (.A1(net242),
    .A2(net237),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06714_ (.I(_01044_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06715_ (.A1(_01605_),
    .A2(_01501_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06716_ (.A1(_01640_),
    .A2(_01348_),
    .B(_01641_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06717_ (.I(_01642_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06718_ (.A1(_01604_),
    .A2(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06719_ (.A1(_01639_),
    .A2(_01644_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06720_ (.A1(_01638_),
    .A2(_01645_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06721_ (.A1(net249),
    .A2(_01617_),
    .B(_01600_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06722_ (.A1(_01637_),
    .A2(_01627_),
    .B1(_01646_),
    .B2(_01647_),
    .ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06723_ (.I(_01388_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06724_ (.A1(net243),
    .A2(_01602_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06725_ (.A1(_01640_),
    .A2(_01031_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06726_ (.A1(_01640_),
    .A2(net347),
    .B(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06727_ (.A1(_01544_),
    .A2(_01651_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06728_ (.A1(_01649_),
    .A2(_01652_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06729_ (.A1(net250),
    .A2(_01078_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06730_ (.A1(_01551_),
    .A2(_01653_),
    .B(_01654_),
    .C(_01612_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06731_ (.A1(_01648_),
    .A2(_01601_),
    .B(_01655_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06732_ (.I(_00805_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06733_ (.I(_01656_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06734_ (.A1(net244),
    .A2(_01007_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06735_ (.A1(_01640_),
    .A2(_01026_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06736_ (.A1(_01606_),
    .A2(_00805_),
    .B(_01659_),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06737_ (.A1(_01543_),
    .A2(_01660_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06738_ (.A1(_01658_),
    .A2(_01661_),
    .B(_01527_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06739_ (.A1(net251),
    .A2(_01617_),
    .B(_01531_),
    .C(_01662_),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06740_ (.A1(_01657_),
    .A2(_01601_),
    .B(_01663_),
    .ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06741_ (.I(_01418_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06742_ (.A1(net245),
    .A2(_01602_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06743_ (.I(_00662_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06744_ (.I(_00764_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06745_ (.A1(_01666_),
    .A2(_01419_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06746_ (.A1(_01666_),
    .A2(_01667_),
    .B(_01668_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06747_ (.A1(_01604_),
    .A2(_01669_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06748_ (.A1(_01665_),
    .A2(_01670_),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06749_ (.A1(_01638_),
    .A2(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06750_ (.A1(net252),
    .A2(_01617_),
    .B(_01600_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06751_ (.A1(_01664_),
    .A2(_01627_),
    .B1(_01672_),
    .B2(_01673_),
    .ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06752_ (.I(_00738_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06753_ (.A1(net246),
    .A2(_01007_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06754_ (.A1(_01666_),
    .A2(_00935_),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06755_ (.A1(_01666_),
    .A2(_00727_),
    .B(_01676_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06756_ (.A1(_01543_),
    .A2(_01677_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06757_ (.A1(_01675_),
    .A2(_01678_),
    .B(_01078_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06758_ (.A1(net253),
    .A2(_01527_),
    .B(_01531_),
    .C(_01679_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06759_ (.A1(_01674_),
    .A2(_01627_),
    .B(_01680_),
    .ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06760_ (.I(\as2650.debug_psu[2] ),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06761_ (.I(_01681_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06762_ (.I(\as2650.debug_psu[3] ),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06763_ (.A1(_01682_),
    .A2(_01683_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06764_ (.I(_01684_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06765_ (.A1(\as2650.debug_psu[0] ),
    .A2(\as2650.debug_psu[1] ),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06766_ (.I(_01686_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06767_ (.I(_01687_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06768_ (.I(_01688_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06769_ (.I(_01689_),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06770_ (.I(_01690_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06771_ (.I(_01691_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06772_ (.I(_01692_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06773_ (.I(_01693_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06774_ (.I(_01236_),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06775_ (.A1(_01695_),
    .A2(_01100_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06776_ (.I(_01696_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06777_ (.A1(_01196_),
    .A2(_01164_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06778_ (.A1(_01698_),
    .A2(_01284_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06779_ (.A1(_01509_),
    .A2(_01699_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06780_ (.I(_01700_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06781_ (.I(_01302_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06782_ (.I(_01163_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06783_ (.A1(_01278_),
    .A2(_01703_),
    .A3(_01364_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06784_ (.A1(_01171_),
    .A2(_01704_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06785_ (.A1(_01250_),
    .A2(_01702_),
    .A3(_01705_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06786_ (.I(_01706_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06787_ (.A1(_01253_),
    .A2(_01455_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06788_ (.A1(_01262_),
    .A2(_01238_),
    .A3(_01323_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06789_ (.A1(_01704_),
    .A2(_01709_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06790_ (.A1(_01505_),
    .A2(_01707_),
    .B1(_01708_),
    .B2(_01710_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06791_ (.A1(_01697_),
    .A2(_01701_),
    .B(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06792_ (.I(_01712_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06793_ (.A1(_01685_),
    .A2(_01694_),
    .A3(_01713_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06794_ (.I(_01714_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06795_ (.I(_01715_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06796_ (.I(_01711_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06797_ (.I(_01717_),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06798_ (.I(\as2650.PC[0] ),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06799_ (.I(_01719_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06800_ (.I(_01720_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06801_ (.I(_00645_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06802_ (.I(\as2650.is_interrupt_cycle ),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06803_ (.A1(_01722_),
    .A2(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06804_ (.I(_01724_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06805_ (.A1(_01721_),
    .A2(_01725_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06806_ (.I(_01131_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06807_ (.A1(_01082_),
    .A2(_01573_),
    .ZN(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06808_ (.I(_01728_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06809_ (.A1(_01727_),
    .A2(_01509_),
    .A3(_01699_),
    .A4(_01729_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06810_ (.I(_01730_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06811_ (.I(_01730_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06812_ (.A1(net188),
    .A2(_01732_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06813_ (.I(_01711_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06814_ (.A1(_01558_),
    .A2(_01731_),
    .B(_01733_),
    .C(_01734_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06815_ (.A1(_01718_),
    .A2(_01726_),
    .B(_01735_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06816_ (.I(_01736_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06817_ (.I(_01714_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06818_ (.I(_01738_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06819_ (.A1(\as2650.stack[12][0] ),
    .A2(_01739_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06820_ (.A1(_01716_),
    .A2(_01737_),
    .B(_01740_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06821_ (.I(_01725_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06822_ (.I(_01724_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06823_ (.A1(\as2650.PC[0] ),
    .A2(\as2650.PC[1] ),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06824_ (.I(_01743_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06825_ (.A1(_01742_),
    .A2(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06826_ (.A1(_00606_),
    .A2(_01741_),
    .B(_01745_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06827_ (.I(_00872_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06828_ (.I(_01204_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06829_ (.I(_01748_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06830_ (.I(_01696_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06831_ (.A1(_01749_),
    .A2(_01750_),
    .A3(_01700_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06832_ (.I(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06833_ (.I(_01752_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06834_ (.I(\as2650.debug_psl[1] ),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06835_ (.I(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06836_ (.I(_01751_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06837_ (.A1(_01755_),
    .A2(_01756_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06838_ (.A1(_01747_),
    .A2(_01753_),
    .B(_01757_),
    .C(_01734_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06839_ (.A1(_01718_),
    .A2(_01746_),
    .B(_01758_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06840_ (.I(_01759_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06841_ (.A1(\as2650.stack[12][1] ),
    .A2(_01739_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06842_ (.A1(_01716_),
    .A2(_01760_),
    .B(_01761_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06843_ (.I(\as2650.PC[1] ),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06844_ (.A1(_01719_),
    .A2(_01762_),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06845_ (.A1(_00610_),
    .A2(_01763_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06846_ (.I(_01764_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06847_ (.A1(_01742_),
    .A2(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06848_ (.A1(_00610_),
    .A2(_01741_),
    .B(_01766_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06849_ (.I(_00895_),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06850_ (.I(_01768_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06851_ (.I(_01752_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06852_ (.I(\as2650.debug_psl[2] ),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06853_ (.I(_01771_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06854_ (.I(_01751_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06855_ (.A1(_01772_),
    .A2(_01773_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06856_ (.A1(_01769_),
    .A2(_01770_),
    .B(_01774_),
    .C(_01717_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06857_ (.A1(_01718_),
    .A2(_01767_),
    .B(_01775_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06858_ (.I(_01776_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06859_ (.A1(\as2650.stack[12][2] ),
    .A2(_01739_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06860_ (.A1(_01716_),
    .A2(_01777_),
    .B(_01778_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06861_ (.I(\as2650.debug_psl[3] ),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _06862_ (.I(_01779_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06863_ (.A1(net214),
    .A2(_01732_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06864_ (.I(_01711_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06865_ (.I(_01782_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06866_ (.A1(_01780_),
    .A2(_01731_),
    .B(_01781_),
    .C(_01783_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06867_ (.A1(_01722_),
    .A2(_01723_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06868_ (.I(_01785_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06869_ (.I(_01786_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06870_ (.I(\as2650.PC[3] ),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06871_ (.I(\as2650.PC[2] ),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06872_ (.A1(_01719_),
    .A2(_01762_),
    .A3(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06873_ (.A1(_01788_),
    .A2(_01790_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06874_ (.I(_01791_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06875_ (.I(_01785_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06876_ (.A1(_01788_),
    .A2(_01793_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06877_ (.A1(_01238_),
    .A2(_01243_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06878_ (.A1(_01708_),
    .A2(_01710_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06879_ (.A1(_01795_),
    .A2(_01706_),
    .B(_01796_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06880_ (.I(_01797_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06881_ (.A1(_01787_),
    .A2(_01792_),
    .B(_01794_),
    .C(_01798_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06882_ (.A1(_01784_),
    .A2(_01799_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06883_ (.I(_01800_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06884_ (.A1(\as2650.stack[12][3] ),
    .A2(_01739_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06885_ (.A1(_01716_),
    .A2(_01801_),
    .B(_01802_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06886_ (.I(_01715_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06887_ (.I(_00923_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06888_ (.I(_01752_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06889_ (.I(_00694_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06890_ (.I(_01806_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06891_ (.I(_01807_),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06892_ (.I(_01752_),
    .Z(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06893_ (.A1(_01808_),
    .A2(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06894_ (.A1(_01804_),
    .A2(_01805_),
    .B(_01810_),
    .C(_01783_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06895_ (.I(\as2650.PC[4] ),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06896_ (.I(_01812_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06897_ (.A1(_00602_),
    .A2(_01790_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06898_ (.A1(_01812_),
    .A2(_01814_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06899_ (.I(_01815_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06900_ (.A1(_01725_),
    .A2(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06901_ (.A1(_01813_),
    .A2(_01741_),
    .B(_01817_),
    .C(_01798_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06902_ (.A1(_01811_),
    .A2(_01818_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06903_ (.I(_01819_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06904_ (.I(_01738_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06905_ (.A1(\as2650.stack[12][4] ),
    .A2(_01821_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06906_ (.A1(_01803_),
    .A2(_01820_),
    .B(_01822_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06907_ (.I(_00803_),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06908_ (.A1(_01569_),
    .A2(_01809_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06909_ (.A1(_01823_),
    .A2(_01805_),
    .B(_01824_),
    .C(_01783_),
    .ZN(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06910_ (.I(\as2650.PC[5] ),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06911_ (.A1(\as2650.PC[4] ),
    .A2(_01826_),
    .A3(_01814_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06912_ (.A1(_01812_),
    .A2(_01814_),
    .B(_01826_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06913_ (.A1(_01827_),
    .A2(_01828_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06914_ (.I(_01829_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06915_ (.I(_01826_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06916_ (.A1(_01831_),
    .A2(_01793_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06917_ (.A1(_01787_),
    .A2(_01830_),
    .B(_01832_),
    .C(_01798_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06918_ (.A1(_01825_),
    .A2(_01833_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06919_ (.I(_01834_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06920_ (.A1(\as2650.stack[12][5] ),
    .A2(_01821_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06921_ (.A1(_01803_),
    .A2(_01835_),
    .B(_01836_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06922_ (.I(_01667_),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06923_ (.I(_01837_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06924_ (.A1(_01560_),
    .A2(_01809_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06925_ (.I(_01782_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06926_ (.A1(_01838_),
    .A2(_01805_),
    .B(_01839_),
    .C(_01840_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06927_ (.I(_01797_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06928_ (.I(_01842_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06929_ (.I(\as2650.PC[6] ),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06930_ (.A1(_01844_),
    .A2(_01827_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06931_ (.I(_01845_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06932_ (.A1(_01742_),
    .A2(_01846_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06933_ (.I(_01844_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06934_ (.I(_01786_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06935_ (.A1(_01848_),
    .A2(_01849_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06936_ (.A1(_01843_),
    .A2(_01847_),
    .A3(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06937_ (.A1(_01841_),
    .A2(_01851_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06938_ (.I(_01852_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06939_ (.A1(\as2650.stack[12][6] ),
    .A2(_01821_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06940_ (.A1(_01803_),
    .A2(_01853_),
    .B(_01854_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06941_ (.I(_00727_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06942_ (.I(_01855_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06943_ (.I(_01856_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06944_ (.A1(_01565_),
    .A2(_01809_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06945_ (.A1(_01857_),
    .A2(_01805_),
    .B(_01858_),
    .C(_01840_),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06946_ (.I(\as2650.PC[7] ),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06947_ (.A1(_01844_),
    .A2(_01860_),
    .A3(_01827_),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06948_ (.I(_01861_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06949_ (.A1(_01844_),
    .A2(_01827_),
    .B(_01860_),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06950_ (.A1(_01862_),
    .A2(_01863_),
    .Z(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06951_ (.I(_01864_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06952_ (.A1(_01860_),
    .A2(_01793_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06953_ (.A1(_01787_),
    .A2(_01865_),
    .B(_01866_),
    .C(_01798_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06954_ (.A1(_01859_),
    .A2(_01867_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06955_ (.I(_01868_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06956_ (.A1(\as2650.stack[12][7] ),
    .A2(_01821_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06957_ (.A1(_01803_),
    .A2(_01869_),
    .B(_01870_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06958_ (.I(_01715_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06959_ (.I(\as2650.debug_psu[0] ),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06960_ (.I(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06961_ (.I(_01873_),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06962_ (.A1(net219),
    .A2(_01732_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06963_ (.A1(_01874_),
    .A2(_01731_),
    .B(_01875_),
    .C(_01840_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06964_ (.I(\as2650.PC[8] ),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06965_ (.A1(_01877_),
    .A2(_01862_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06966_ (.I(_01877_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06967_ (.A1(_01879_),
    .A2(_01793_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06968_ (.A1(_01787_),
    .A2(_01878_),
    .B(_01880_),
    .C(_01842_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06969_ (.A1(_01876_),
    .A2(_01881_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06970_ (.I(_01882_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06971_ (.I(_01738_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06972_ (.A1(\as2650.stack[12][8] ),
    .A2(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06973_ (.A1(_01871_),
    .A2(_01883_),
    .B(_01885_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06974_ (.I(\as2650.debug_psu[1] ),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06975_ (.I(_01886_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06976_ (.A1(_01887_),
    .A2(_01756_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06977_ (.A1(_01351_),
    .A2(_01753_),
    .B(_01888_),
    .C(_01840_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06978_ (.I(\as2650.PC[9] ),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06979_ (.A1(\as2650.PC[8] ),
    .A2(_01862_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06980_ (.A1(_01890_),
    .A2(_01891_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06981_ (.I(_01892_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06982_ (.A1(_01742_),
    .A2(_01893_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06983_ (.I(_01890_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06984_ (.A1(_01895_),
    .A2(_01849_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06985_ (.A1(_01843_),
    .A2(_01894_),
    .A3(_01896_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06986_ (.A1(_01889_),
    .A2(_01897_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06987_ (.I(_01898_),
    .Z(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06988_ (.A1(\as2650.stack[12][9] ),
    .A2(_01884_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06989_ (.A1(_01871_),
    .A2(_01899_),
    .B(_01900_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06990_ (.I(_01682_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06991_ (.I(_01901_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06992_ (.A1(_01902_),
    .A2(_01756_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06993_ (.A1(_01369_),
    .A2(_01753_),
    .B(_01903_),
    .C(_01734_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06994_ (.I(\as2650.PC[10] ),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06995_ (.A1(\as2650.PC[8] ),
    .A2(_01890_),
    .A3(_01861_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06996_ (.A1(_01905_),
    .A2(_01906_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06997_ (.I(_01907_),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06998_ (.I(_01908_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06999_ (.A1(_01905_),
    .A2(_01786_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07000_ (.A1(_01849_),
    .A2(_01909_),
    .B(_01910_),
    .C(_01842_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07001_ (.A1(_01904_),
    .A2(_01911_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07002_ (.I(_01912_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07003_ (.A1(\as2650.stack[12][10] ),
    .A2(_01884_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07004_ (.A1(_01871_),
    .A2(_01913_),
    .B(_01914_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07005_ (.I(\as2650.PC[11] ),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07006_ (.I(_01915_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07007_ (.I(_01905_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07008_ (.A1(_01917_),
    .A2(_01906_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07009_ (.A1(_01915_),
    .A2(_01918_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07010_ (.I(_01919_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07011_ (.A1(_01725_),
    .A2(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07012_ (.A1(_01916_),
    .A2(_01741_),
    .B(_01921_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07013_ (.I(_01683_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07014_ (.I(_01923_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07015_ (.A1(net190),
    .A2(_01732_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07016_ (.A1(_01924_),
    .A2(_01731_),
    .B(_01925_),
    .C(_01717_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07017_ (.A1(_01783_),
    .A2(_01922_),
    .B(_01926_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07018_ (.I(_01927_),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07019_ (.A1(\as2650.stack[12][11] ),
    .A2(_01884_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07020_ (.A1(_01871_),
    .A2(_01928_),
    .B(_01929_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07021_ (.I(_01715_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07022_ (.I(\as2650.debug_psu[4] ),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07023_ (.A1(_01931_),
    .A2(_01756_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07024_ (.A1(_00915_),
    .A2(_01753_),
    .B(_01932_),
    .C(_01734_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07025_ (.I(\as2650.PC[12] ),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07026_ (.A1(_01915_),
    .A2(_01918_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _07027_ (.A1(_01934_),
    .A2(_01935_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07028_ (.A1(_01934_),
    .A2(_01786_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07029_ (.A1(_01849_),
    .A2(_01936_),
    .B(_01937_),
    .C(_01842_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07030_ (.A1(_01933_),
    .A2(_01938_),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07031_ (.I(_01939_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07032_ (.I(_01738_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07033_ (.A1(\as2650.stack[12][12] ),
    .A2(_01941_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07034_ (.A1(_01930_),
    .A2(_01940_),
    .B(_01942_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _07035_ (.I(_01092_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07036_ (.A1(net192),
    .A2(_01773_),
    .B(_01782_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07037_ (.A1(_01943_),
    .A2(_01770_),
    .B(_01944_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07038_ (.A1(_00958_),
    .A2(_01843_),
    .B(_01945_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07039_ (.I(_01946_),
    .Z(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07040_ (.A1(\as2650.stack[12][13] ),
    .A2(_01941_),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07041_ (.A1(_01930_),
    .A2(_01947_),
    .B(_01948_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07042_ (.I(\as2650.page_reg[1] ),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _07043_ (.I(net306),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07044_ (.A1(net193),
    .A2(_01773_),
    .B(_01782_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07045_ (.A1(_01950_),
    .A2(_01770_),
    .B(_01951_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07046_ (.A1(_01949_),
    .A2(_01843_),
    .B(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07047_ (.I(_01953_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07048_ (.A1(\as2650.stack[12][14] ),
    .A2(_01941_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07049_ (.A1(_01930_),
    .A2(_01954_),
    .B(_01955_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07050_ (.A1(\as2650.debug_psu[7] ),
    .A2(_01773_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07051_ (.A1(_00722_),
    .A2(_01770_),
    .B(_01956_),
    .C(_01717_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07052_ (.A1(\as2650.page_reg[2] ),
    .A2(_01718_),
    .B(_01957_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07053_ (.I(_01958_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07054_ (.A1(\as2650.stack[12][15] ),
    .A2(_01941_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07055_ (.A1(_01930_),
    .A2(_01959_),
    .B(_01960_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07056_ (.I(_01712_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07057_ (.A1(_01901_),
    .A2(_01924_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07058_ (.A1(_01872_),
    .A2(_01886_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07059_ (.I(_01963_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07060_ (.I(_01964_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07061_ (.I(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07062_ (.I(_01966_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07063_ (.I(_01967_),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07064_ (.I(_01968_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07065_ (.I(_01969_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07066_ (.A1(_01961_),
    .A2(_01962_),
    .A3(_01970_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07067_ (.I(_01971_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07068_ (.I(_01972_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07069_ (.I(_01971_),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07070_ (.I(_01974_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07071_ (.A1(\as2650.stack[11][0] ),
    .A2(_01975_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07072_ (.A1(_01737_),
    .A2(_01973_),
    .B(_01976_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07073_ (.A1(\as2650.stack[11][1] ),
    .A2(_01975_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07074_ (.A1(_01760_),
    .A2(_01973_),
    .B(_01977_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07075_ (.A1(\as2650.stack[11][2] ),
    .A2(_01975_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07076_ (.A1(_01777_),
    .A2(_01973_),
    .B(_01978_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07077_ (.A1(\as2650.stack[11][3] ),
    .A2(_01975_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07078_ (.A1(_01801_),
    .A2(_01973_),
    .B(_01979_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07079_ (.I(_01972_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07080_ (.I(_01974_),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07081_ (.A1(\as2650.stack[11][4] ),
    .A2(_01981_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07082_ (.A1(_01820_),
    .A2(_01980_),
    .B(_01982_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07083_ (.A1(\as2650.stack[11][5] ),
    .A2(_01981_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07084_ (.A1(_01835_),
    .A2(_01980_),
    .B(_01983_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07085_ (.A1(\as2650.stack[11][6] ),
    .A2(_01981_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07086_ (.A1(_01853_),
    .A2(_01980_),
    .B(_01984_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07087_ (.A1(\as2650.stack[11][7] ),
    .A2(_01981_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07088_ (.A1(_01869_),
    .A2(_01980_),
    .B(_01985_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07089_ (.I(_01972_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07090_ (.I(_01974_),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07091_ (.A1(\as2650.stack[11][8] ),
    .A2(_01987_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07092_ (.A1(_01883_),
    .A2(_01986_),
    .B(_01988_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07093_ (.A1(\as2650.stack[11][9] ),
    .A2(_01987_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07094_ (.A1(_01899_),
    .A2(_01986_),
    .B(_01989_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07095_ (.A1(\as2650.stack[11][10] ),
    .A2(_01987_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07096_ (.A1(_01913_),
    .A2(_01986_),
    .B(_01990_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07097_ (.A1(\as2650.stack[11][11] ),
    .A2(_01987_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07098_ (.A1(_01928_),
    .A2(_01986_),
    .B(_01991_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07099_ (.I(_01972_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07100_ (.I(_01974_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07101_ (.A1(\as2650.stack[11][12] ),
    .A2(_01993_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07102_ (.A1(_01940_),
    .A2(_01992_),
    .B(_01994_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07103_ (.A1(\as2650.stack[11][13] ),
    .A2(_01993_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07104_ (.A1(_01947_),
    .A2(_01992_),
    .B(_01995_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07105_ (.A1(\as2650.stack[11][14] ),
    .A2(_01993_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07106_ (.A1(_01954_),
    .A2(_01992_),
    .B(_01996_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07107_ (.A1(\as2650.stack[11][15] ),
    .A2(_01993_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07108_ (.A1(_01959_),
    .A2(_01992_),
    .B(_01997_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07109_ (.I(_01307_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07110_ (.A1(_01998_),
    .A2(_01266_),
    .A3(_01469_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07111_ (.I(_01472_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07112_ (.I(_02000_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07113_ (.A1(_01181_),
    .A2(_01324_),
    .A3(_01454_),
    .A4(_02001_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07114_ (.I(_01086_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07115_ (.I(_02003_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07116_ (.A1(_01999_),
    .A2(_02002_),
    .B(_02004_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07117_ (.A1(net104),
    .A2(net71),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07118_ (.A1(wb_feedback_delay),
    .A2(_02005_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07119_ (.A1(net105),
    .A2(_02006_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07120_ (.A1(net70),
    .A2(_02007_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07121_ (.I(net69),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07122_ (.I(net68),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07123_ (.A1(_02009_),
    .A2(_02010_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07124_ (.A1(net66),
    .A2(net67),
    .A3(_02011_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07125_ (.A1(_02008_),
    .A2(_02012_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07126_ (.I(_02013_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07127_ (.I(_02014_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07128_ (.I0(net72),
    .I1(net122),
    .S(_02015_),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07129_ (.I(_02016_),
    .Z(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07130_ (.I0(net83),
    .I1(net129),
    .S(_02015_),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07131_ (.I(_02017_),
    .Z(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07132_ (.I0(net94),
    .I1(net130),
    .S(_02015_),
    .Z(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07133_ (.I(_02018_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07134_ (.I0(net97),
    .I1(net131),
    .S(_02015_),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07135_ (.I(_02019_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07136_ (.I(_02014_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07137_ (.I0(net98),
    .I1(net132),
    .S(_02020_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07138_ (.I(_02021_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07139_ (.I0(net99),
    .I1(net133),
    .S(_02020_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07140_ (.I(_02022_),
    .Z(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07141_ (.I0(net100),
    .I1(net134),
    .S(_02020_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07142_ (.I(_02023_),
    .Z(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07143_ (.I0(net101),
    .I1(net135),
    .S(_02020_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07144_ (.I(_02024_),
    .Z(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07145_ (.I(_02014_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07146_ (.I0(net102),
    .I1(net136),
    .S(_02025_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07147_ (.I(_02026_),
    .Z(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07148_ (.I0(net103),
    .I1(net137),
    .S(_02025_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07149_ (.I(_02027_),
    .Z(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07150_ (.I0(net73),
    .I1(net123),
    .S(_02025_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07151_ (.I(net409),
    .Z(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07152_ (.I0(net74),
    .I1(net124),
    .S(_02025_),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07153_ (.I(_02029_),
    .Z(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07154_ (.I(_02014_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07155_ (.I0(net75),
    .I1(net125),
    .S(_02030_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07156_ (.I(_02031_),
    .Z(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07157_ (.I0(net76),
    .I1(net126),
    .S(_02030_),
    .Z(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07158_ (.I(_02032_),
    .Z(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07159_ (.I0(net77),
    .I1(net127),
    .S(_02030_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07160_ (.I(_02033_),
    .Z(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07161_ (.I0(net78),
    .I1(net128),
    .S(_02030_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07162_ (.I(_02034_),
    .Z(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07163_ (.I(_02013_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07164_ (.I(_02035_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07165_ (.I0(net79),
    .I1(net106),
    .S(_02036_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07166_ (.I(_02037_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07167_ (.I0(net80),
    .I1(net113),
    .S(_02036_),
    .Z(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07168_ (.I(_02038_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07169_ (.I0(net81),
    .I1(net114),
    .S(_02036_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07170_ (.I(_02039_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07171_ (.I0(net82),
    .I1(net115),
    .S(_02036_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07172_ (.I(_02040_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07173_ (.I(_02035_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07174_ (.I0(net84),
    .I1(net116),
    .S(_02041_),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07175_ (.I(_02042_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07176_ (.I0(net85),
    .I1(net117),
    .S(_02041_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07177_ (.I(_02043_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07178_ (.I0(net86),
    .I1(net118),
    .S(_02041_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07179_ (.I(_02044_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07180_ (.I0(net87),
    .I1(net119),
    .S(_02041_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07181_ (.I(_02045_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07182_ (.I(_02035_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07183_ (.I0(net88),
    .I1(net120),
    .S(_02046_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07184_ (.I(_02047_),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07185_ (.I0(net89),
    .I1(net121),
    .S(_02046_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07186_ (.I(_02048_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07187_ (.I0(net90),
    .I1(net107),
    .S(_02046_),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07188_ (.I(_02049_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07189_ (.I0(net91),
    .I1(net108),
    .S(_02046_),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07190_ (.I(_02050_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07191_ (.I(_02035_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07192_ (.I0(net92),
    .I1(net109),
    .S(_02051_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07193_ (.I(_02052_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07194_ (.I0(net93),
    .I1(net110),
    .S(_02051_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07195_ (.I(_02053_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07196_ (.I0(net95),
    .I1(net111),
    .S(_02051_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07197_ (.I(_02054_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07198_ (.I0(net96),
    .I1(net112),
    .S(_02051_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07199_ (.I(_02055_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07200_ (.I(net69),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07201_ (.A1(_02056_),
    .A2(_02008_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07202_ (.I(_02057_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07203_ (.I(_02058_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07204_ (.I(_02058_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07205_ (.A1(net102),
    .A2(_02060_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07206_ (.I(net66),
    .Z(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07207_ (.I(_02062_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07208_ (.A1(_01119_),
    .A2(_02059_),
    .B(_02061_),
    .C(_02063_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07209_ (.I(net67),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07210_ (.A1(net105),
    .A2(_02006_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07211_ (.I(net70),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07212_ (.A1(_02056_),
    .A2(_02066_),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07213_ (.A1(_02010_),
    .A2(_02064_),
    .A3(_02065_),
    .A4(_02067_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07214_ (.A1(_02062_),
    .A2(_02068_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07215_ (.I0(net159),
    .I1(net72),
    .S(_02069_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07216_ (.I(_02070_),
    .Z(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07217_ (.I0(net160),
    .I1(net83),
    .S(_02069_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07218_ (.I(_02071_),
    .Z(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07219_ (.I0(net161),
    .I1(net94),
    .S(_02069_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07220_ (.I(_02072_),
    .Z(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07221_ (.I(net66),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07222_ (.I(_02073_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07223_ (.I(_02074_),
    .Z(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07224_ (.A1(_02075_),
    .A2(wb_feedback_delay),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07225_ (.I(_02076_),
    .Z(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07226_ (.A1(wb_feedback_delay),
    .A2(net105),
    .A3(_02005_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07227_ (.I(_02077_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07228_ (.I(_02078_),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07229_ (.I(_02079_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07230_ (.I(_02066_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07231_ (.I(_02081_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07232_ (.I(_02056_),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07233_ (.I(_02064_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07234_ (.A1(_02084_),
    .A2(net159),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07235_ (.I(net67),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07236_ (.I(_02011_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07237_ (.A1(_02086_),
    .A2(net122),
    .B(_02087_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07238_ (.A1(_01561_),
    .A2(_02083_),
    .B1(_02085_),
    .B2(_02088_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07239_ (.I(_02066_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07240_ (.I(\wb_counter[0] ),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07241_ (.A1(_02090_),
    .A2(_02091_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07242_ (.A1(_02082_),
    .A2(_02089_),
    .B(_02092_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07243_ (.I(_02077_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07244_ (.I(_02094_),
    .Z(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07245_ (.A1(net266),
    .A2(_02095_),
    .B(_02075_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07246_ (.A1(_02080_),
    .A2(_02093_),
    .B(_02096_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07247_ (.I(wb_debug_carry),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07248_ (.A1(_02084_),
    .A2(net160),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07249_ (.A1(_02086_),
    .A2(net129),
    .B(_02087_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07250_ (.A1(_02097_),
    .A2(_02083_),
    .B1(_02098_),
    .B2(_02099_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07251_ (.I(\wb_counter[1] ),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07252_ (.A1(_02090_),
    .A2(_02101_),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07253_ (.A1(_02082_),
    .A2(_02100_),
    .B(_02102_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07254_ (.A1(net277),
    .A2(_02095_),
    .B(_02075_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07255_ (.A1(_02080_),
    .A2(_02103_),
    .B(_02104_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07256_ (.A1(_02084_),
    .A2(net161),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07257_ (.A1(_02086_),
    .A2(net130),
    .B(_02087_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07258_ (.A1(_01553_),
    .A2(_02083_),
    .B1(_02105_),
    .B2(_02106_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07259_ (.I(\wb_counter[2] ),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07260_ (.A1(_02090_),
    .A2(_02108_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07261_ (.A1(_02082_),
    .A2(_02107_),
    .B(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07262_ (.A1(net288),
    .A2(_02095_),
    .B(_02075_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07263_ (.A1(_02080_),
    .A2(_02110_),
    .B(_02111_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07264_ (.I(net70),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07265_ (.I(_02112_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07266_ (.I(_02113_),
    .Z(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07267_ (.I(_02112_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07268_ (.I(_02115_),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07269_ (.A1(_02010_),
    .A2(_02086_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07270_ (.I(_02117_),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07271_ (.I(_02118_),
    .Z(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07272_ (.A1(net68),
    .A2(net67),
    .B(net69),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07273_ (.I(_02120_),
    .Z(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07274_ (.I(_02121_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07275_ (.A1(net131),
    .A2(_02119_),
    .B(_02122_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07276_ (.I(_02056_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07277_ (.A1(\web_behavior[1] ),
    .A2(_02124_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07278_ (.A1(_02116_),
    .A2(_02123_),
    .A3(_02125_),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07279_ (.A1(_02114_),
    .A2(\wb_counter[3] ),
    .B(_02126_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07280_ (.I(_02074_),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07281_ (.A1(net291),
    .A2(_02095_),
    .B(_02128_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07282_ (.A1(_02080_),
    .A2(_02127_),
    .B(_02129_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07283_ (.I(_02079_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07284_ (.I(\wb_counter[4] ),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07285_ (.A1(net132),
    .A2(_02119_),
    .B(_02122_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07286_ (.A1(wb_reset_override_en),
    .A2(_02124_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07287_ (.A1(_02116_),
    .A2(_02132_),
    .A3(_02133_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07288_ (.A1(_02114_),
    .A2(_02131_),
    .B(_02134_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07289_ (.I(_02077_),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07290_ (.I(_02136_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07291_ (.A1(net292),
    .A2(_02137_),
    .B(_02128_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07292_ (.A1(_02130_),
    .A2(_02135_),
    .B(_02138_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07293_ (.I(_02118_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07294_ (.A1(net133),
    .A2(_02139_),
    .B(_02122_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07295_ (.I(net69),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07296_ (.A1(wb_reset_override),
    .A2(_02141_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07297_ (.A1(_02116_),
    .A2(_02140_),
    .A3(_02142_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07298_ (.A1(_02114_),
    .A2(\wb_counter[5] ),
    .B(_02143_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07299_ (.A1(net293),
    .A2(_02137_),
    .B(_02128_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07300_ (.A1(_02130_),
    .A2(_02144_),
    .B(_02145_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07301_ (.I(_02009_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07302_ (.I(_02146_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07303_ (.I(_02112_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07304_ (.I(_02118_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07305_ (.I(_02121_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07306_ (.A1(net134),
    .A2(_02149_),
    .B(_02150_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07307_ (.A1(net165),
    .A2(_02147_),
    .B(_02148_),
    .C(_02151_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07308_ (.A1(_02114_),
    .A2(\wb_counter[6] ),
    .B(_02152_),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07309_ (.A1(net294),
    .A2(_02137_),
    .B(_02128_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07310_ (.A1(_02130_),
    .A2(_02153_),
    .B(_02154_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07311_ (.I(_02113_),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07312_ (.A1(net135),
    .A2(_02139_),
    .B(_02122_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07313_ (.A1(net182),
    .A2(_02141_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07314_ (.A1(_02116_),
    .A2(_02156_),
    .A3(_02157_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07315_ (.A1(_02155_),
    .A2(\wb_counter[7] ),
    .B(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07316_ (.I(_02074_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07317_ (.A1(net295),
    .A2(_02137_),
    .B(_02160_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07318_ (.A1(_02130_),
    .A2(_02159_),
    .B(_02161_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07319_ (.I(_02079_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07320_ (.A1(net136),
    .A2(_02149_),
    .B(_02150_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07321_ (.A1(_01119_),
    .A2(_02147_),
    .B(_02148_),
    .C(_02163_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07322_ (.A1(_02155_),
    .A2(\wb_counter[8] ),
    .B(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07323_ (.I(_02136_),
    .Z(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07324_ (.A1(net296),
    .A2(_02166_),
    .B(_02160_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07325_ (.A1(_02162_),
    .A2(_02165_),
    .B(_02167_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07326_ (.I(_02117_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07327_ (.A1(net137),
    .A2(_02168_),
    .B(_02150_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07328_ (.I(_02112_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07329_ (.A1(_02147_),
    .A2(_01558_),
    .B(_02169_),
    .C(_02170_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07330_ (.A1(_02155_),
    .A2(\wb_counter[9] ),
    .B(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07331_ (.A1(net297),
    .A2(_02166_),
    .B(_02160_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07332_ (.A1(_02162_),
    .A2(_02172_),
    .B(_02173_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07333_ (.I(_02115_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07334_ (.I(_02121_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07335_ (.A1(net123),
    .A2(_02139_),
    .B(_02175_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07336_ (.A1(_02083_),
    .A2(_01755_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07337_ (.A1(_02174_),
    .A2(_02176_),
    .A3(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07338_ (.A1(_02155_),
    .A2(\wb_counter[10] ),
    .B(_02178_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07339_ (.A1(net267),
    .A2(_02166_),
    .B(_02160_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07340_ (.A1(_02162_),
    .A2(_02179_),
    .B(_02180_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07341_ (.I(_02113_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07342_ (.A1(net124),
    .A2(_02139_),
    .B(_02175_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07343_ (.I(_02141_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07344_ (.A1(_02183_),
    .A2(_01772_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07345_ (.A1(_02174_),
    .A2(_02182_),
    .A3(_02184_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07346_ (.A1(_02181_),
    .A2(\wb_counter[11] ),
    .B(_02185_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07347_ (.I(_02073_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07348_ (.I(_02187_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07349_ (.A1(net268),
    .A2(_02166_),
    .B(_02188_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07350_ (.A1(_02162_),
    .A2(_02186_),
    .B(_02189_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07351_ (.I(_02078_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07352_ (.I(_02190_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07353_ (.I(_02009_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07354_ (.I(_02120_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07355_ (.A1(net125),
    .A2(_02168_),
    .B(_02193_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07356_ (.A1(_02192_),
    .A2(_01780_),
    .B(_02194_),
    .C(_02170_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07357_ (.A1(_02181_),
    .A2(\wb_counter[12] ),
    .B(_02195_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07358_ (.I(_02136_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07359_ (.A1(net269),
    .A2(_02197_),
    .B(_02188_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07360_ (.A1(_02191_),
    .A2(_02196_),
    .B(_02198_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07361_ (.I(_02118_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07362_ (.A1(net126),
    .A2(_02199_),
    .B(_02175_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07363_ (.I(_01808_),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07364_ (.A1(_02201_),
    .A2(_02141_),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07365_ (.A1(_02174_),
    .A2(_02200_),
    .A3(_02202_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07366_ (.A1(_02181_),
    .A2(\wb_counter[13] ),
    .B(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07367_ (.A1(net270),
    .A2(_02197_),
    .B(_02188_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07368_ (.A1(_02191_),
    .A2(_02204_),
    .B(_02205_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07369_ (.A1(net127),
    .A2(_02199_),
    .B(_02175_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07370_ (.A1(_02183_),
    .A2(_01570_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07371_ (.A1(_02174_),
    .A2(_02206_),
    .A3(_02207_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07372_ (.A1(_02181_),
    .A2(\wb_counter[14] ),
    .B(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07373_ (.A1(net271),
    .A2(_02197_),
    .B(_02188_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07374_ (.A1(_02191_),
    .A2(_02209_),
    .B(_02210_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07375_ (.I(_02113_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07376_ (.I(_02115_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07377_ (.I(_02121_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07378_ (.A1(net128),
    .A2(_02199_),
    .B(_02213_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07379_ (.A1(_02183_),
    .A2(_01560_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07380_ (.A1(_02212_),
    .A2(_02214_),
    .A3(_02215_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07381_ (.A1(_02211_),
    .A2(\wb_counter[15] ),
    .B(_02216_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07382_ (.I(_02187_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07383_ (.A1(net272),
    .A2(_02197_),
    .B(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07384_ (.A1(_02191_),
    .A2(_02217_),
    .B(_02219_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07385_ (.I(_02190_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07386_ (.A1(net106),
    .A2(_02199_),
    .B(_02213_),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07387_ (.A1(_02183_),
    .A2(_01565_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07388_ (.A1(_02212_),
    .A2(_02221_),
    .A3(_02222_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07389_ (.A1(_02211_),
    .A2(\wb_counter[16] ),
    .B(_02223_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07390_ (.I(_02136_),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07391_ (.A1(net273),
    .A2(_02225_),
    .B(_02218_),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07392_ (.A1(_02220_),
    .A2(_02224_),
    .B(_02226_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07393_ (.A1(net113),
    .A2(_02168_),
    .B(_02193_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07394_ (.A1(_02192_),
    .A2(_01874_),
    .B(_02227_),
    .C(_02170_),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07395_ (.A1(_02211_),
    .A2(\wb_counter[17] ),
    .B(_02228_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07396_ (.A1(net274),
    .A2(_02225_),
    .B(_02218_),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07397_ (.A1(_02220_),
    .A2(_02229_),
    .B(_02230_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07398_ (.A1(net114),
    .A2(_02149_),
    .B(_02213_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07399_ (.A1(_02124_),
    .A2(_01887_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07400_ (.A1(_02212_),
    .A2(_02231_),
    .A3(_02232_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07401_ (.A1(_02211_),
    .A2(\wb_counter[18] ),
    .B(_02233_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07402_ (.A1(net275),
    .A2(_02225_),
    .B(_02218_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07403_ (.A1(_02220_),
    .A2(_02234_),
    .B(_02235_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07404_ (.I(_02062_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07405_ (.I(_02236_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07406_ (.I(_02077_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07407_ (.I(_02066_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07408_ (.A1(_02084_),
    .A2(net115),
    .A3(_02087_),
    .B1(_01902_),
    .B2(_02146_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07409_ (.A1(_02081_),
    .A2(\wb_counter[19] ),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07410_ (.A1(_02239_),
    .A2(_02240_),
    .B(_02241_),
    .C(_02094_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07411_ (.A1(net276),
    .A2(_02238_),
    .B(_02242_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07412_ (.A1(_02237_),
    .A2(_02243_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07413_ (.I(_02115_),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07414_ (.I(_02117_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07415_ (.A1(net116),
    .A2(_02245_),
    .B(_02193_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07416_ (.A1(_02192_),
    .A2(_01924_),
    .B(_02246_),
    .C(_02170_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07417_ (.A1(_02244_),
    .A2(\wb_counter[20] ),
    .B(_02247_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07418_ (.I(_02187_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07419_ (.A1(net278),
    .A2(_02225_),
    .B(_02249_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07420_ (.A1(_02220_),
    .A2(_02248_),
    .B(_02250_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07421_ (.I(_02190_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07422_ (.A1(net117),
    .A2(_02149_),
    .B(_02213_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07423_ (.A1(_02124_),
    .A2(_01931_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07424_ (.A1(_02212_),
    .A2(_02252_),
    .A3(_02253_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07425_ (.A1(_02244_),
    .A2(\wb_counter[21] ),
    .B(_02254_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07426_ (.I(_02078_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07427_ (.A1(net279),
    .A2(_02256_),
    .B(_02249_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07428_ (.A1(_02251_),
    .A2(_02255_),
    .B(_02257_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07429_ (.A1(net118),
    .A2(_02168_),
    .B(_02150_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07430_ (.A1(_01943_),
    .A2(_02147_),
    .B(_02148_),
    .C(_02258_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07431_ (.A1(_02244_),
    .A2(\wb_counter[22] ),
    .B(_02259_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07432_ (.A1(net280),
    .A2(_02256_),
    .B(_02249_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07433_ (.A1(_02251_),
    .A2(_02260_),
    .B(_02261_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07434_ (.A1(net119),
    .A2(_02245_),
    .B(_02193_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07435_ (.A1(_02192_),
    .A2(_01950_),
    .B(_02262_),
    .C(_02148_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07436_ (.A1(_02244_),
    .A2(\wb_counter[23] ),
    .B(_02263_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07437_ (.A1(net281),
    .A2(_02256_),
    .B(_02249_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07438_ (.A1(_02251_),
    .A2(_02264_),
    .B(_02265_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07439_ (.A1(_02064_),
    .A2(net120),
    .A3(_02011_),
    .B1(\as2650.debug_psu[7] ),
    .B2(_02146_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07440_ (.A1(_02081_),
    .A2(\wb_counter[24] ),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07441_ (.A1(_02239_),
    .A2(_02266_),
    .B(_02267_),
    .C(_02094_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07442_ (.A1(net282),
    .A2(_02238_),
    .B(_02268_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07443_ (.A1(_02237_),
    .A2(_02269_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07444_ (.A1(net121),
    .A2(_02119_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07445_ (.A1(_02010_),
    .A2(_02064_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07446_ (.I(_02067_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07447_ (.A1(_02271_),
    .A2(_02272_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07448_ (.A1(_02082_),
    .A2(\wb_counter[25] ),
    .B1(_02270_),
    .B2(_02273_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07449_ (.I(_02187_),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07450_ (.A1(net283),
    .A2(_02256_),
    .B(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07451_ (.A1(_02251_),
    .A2(_02274_),
    .B(_02276_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07452_ (.I(_02190_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07453_ (.I(_02081_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07454_ (.I(_02245_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07455_ (.A1(net107),
    .A2(_02279_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07456_ (.A1(_02278_),
    .A2(\wb_counter[26] ),
    .B1(_02273_),
    .B2(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07457_ (.I(_02078_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07458_ (.A1(net284),
    .A2(_02282_),
    .B(_02275_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07459_ (.A1(_02277_),
    .A2(_02281_),
    .B(_02283_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07460_ (.A1(net108),
    .A2(_02279_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07461_ (.A1(_02278_),
    .A2(\wb_counter[27] ),
    .B1(_02273_),
    .B2(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07462_ (.A1(net285),
    .A2(_02282_),
    .B(_02275_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07463_ (.A1(_02277_),
    .A2(_02285_),
    .B(_02286_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07464_ (.A1(net109),
    .A2(_02279_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07465_ (.A1(_02278_),
    .A2(\wb_counter[28] ),
    .B1(_02272_),
    .B2(_02287_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07466_ (.A1(net286),
    .A2(_02282_),
    .B(_02275_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07467_ (.A1(_02277_),
    .A2(_02288_),
    .B(_02289_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07468_ (.A1(net110),
    .A2(_02279_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07469_ (.A1(_02278_),
    .A2(\wb_counter[29] ),
    .B1(_02272_),
    .B2(_02290_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07470_ (.I(_02073_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07471_ (.I(_02292_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07472_ (.A1(net287),
    .A2(_02282_),
    .B(_02293_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07473_ (.A1(_02277_),
    .A2(_02291_),
    .B(_02294_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07474_ (.A1(net111),
    .A2(_02119_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07475_ (.A1(_02090_),
    .A2(\wb_counter[30] ),
    .B1(_02273_),
    .B2(_02295_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07476_ (.A1(net289),
    .A2(_02079_),
    .B(_02293_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07477_ (.A1(_02238_),
    .A2(_02296_),
    .B(_02297_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07478_ (.A1(\as2650.wb_hidden_rom_enable ),
    .A2(_02271_),
    .B1(_02245_),
    .B2(net112),
    .C(_02272_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07479_ (.A1(_02239_),
    .A2(\wb_counter[31] ),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07480_ (.A1(_02094_),
    .A2(_02298_),
    .A3(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07481_ (.A1(net290),
    .A2(_02238_),
    .B(_02300_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07482_ (.A1(_02237_),
    .A2(_02301_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07483_ (.A1(_02237_),
    .A2(net427),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07484_ (.A1(net72),
    .A2(_02060_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07485_ (.A1(_01561_),
    .A2(_02059_),
    .B(_02302_),
    .C(_02063_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07486_ (.A1(net83),
    .A2(_02060_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07487_ (.A1(_02097_),
    .A2(_02059_),
    .B(_02303_),
    .C(_02063_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07488_ (.A1(net94),
    .A2(_02058_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07489_ (.A1(_01553_),
    .A2(_02059_),
    .B(_02304_),
    .C(_02063_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07490_ (.I(_02057_),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07491_ (.A1(\web_behavior[1] ),
    .A2(_02305_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07492_ (.A1(_02146_),
    .A2(_02239_),
    .A3(_02007_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07493_ (.A1(net366),
    .A2(_02307_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07494_ (.I(_02062_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07495_ (.A1(_02306_),
    .A2(net367),
    .B(_02309_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07496_ (.A1(wb_reset_override_en),
    .A2(_02305_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07497_ (.A1(net358),
    .A2(_02307_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07498_ (.A1(_02310_),
    .A2(net359),
    .B(_02309_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07499_ (.A1(wb_reset_override),
    .A2(_02305_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07500_ (.A1(net362),
    .A2(_02307_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07501_ (.A1(_02312_),
    .A2(net363),
    .B(_02309_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07502_ (.A1(net100),
    .A2(_02058_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07503_ (.A1(net165),
    .A2(_02305_),
    .B(_02314_),
    .C(_02236_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07504_ (.A1(net182),
    .A2(_02060_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07505_ (.A1(net101),
    .A2(_02307_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07506_ (.A1(_02315_),
    .A2(net370),
    .B(_02309_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07507_ (.I(\as2650.wb_hidden_rom_enable ),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07508_ (.A1(net96),
    .A2(net437),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07509_ (.A1(_02317_),
    .A2(net411),
    .B(_02318_),
    .C(_02236_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07510_ (.A1(net70),
    .A2(_02065_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07511_ (.I(_02319_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07512_ (.I(_02320_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07513_ (.I(_02319_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07514_ (.I(_02322_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07515_ (.A1(net72),
    .A2(_02323_),
    .B(_02293_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07516_ (.A1(\wb_counter[0] ),
    .A2(_02321_),
    .B(_02324_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07517_ (.A1(_02091_),
    .A2(\wb_counter[1] ),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07518_ (.A1(net83),
    .A2(_02323_),
    .B(_02293_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07519_ (.A1(_02321_),
    .A2(_02325_),
    .B(_02326_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07520_ (.A1(\wb_counter[0] ),
    .A2(\wb_counter[1] ),
    .A3(\wb_counter[2] ),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07521_ (.A1(_02091_),
    .A2(_02101_),
    .B(_02108_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07522_ (.A1(_02327_),
    .A2(_02328_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07523_ (.I(_02292_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07524_ (.A1(net94),
    .A2(_02323_),
    .B(_02330_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07525_ (.A1(_02321_),
    .A2(_02329_),
    .B(_02331_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07526_ (.I(_02320_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07527_ (.A1(\wb_counter[3] ),
    .A2(_02327_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07528_ (.A1(net97),
    .A2(_02320_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07529_ (.A1(_02332_),
    .A2(_02333_),
    .B(net433),
    .C(_02236_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07530_ (.I(\wb_counter[3] ),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07531_ (.A1(_02335_),
    .A2(_02327_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07532_ (.A1(_02131_),
    .A2(_02336_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07533_ (.A1(net358),
    .A2(_02323_),
    .B(_02330_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07534_ (.A1(_02321_),
    .A2(_02337_),
    .B(_02338_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07535_ (.I(_02319_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07536_ (.I(_02339_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07537_ (.I(_02340_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07538_ (.A1(_02131_),
    .A2(_02336_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07539_ (.A1(\wb_counter[5] ),
    .A2(_02342_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07540_ (.I(_02322_),
    .Z(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07541_ (.A1(net362),
    .A2(_02344_),
    .B(_02330_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07542_ (.A1(_02341_),
    .A2(_02343_),
    .B(_02345_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07543_ (.A1(_02131_),
    .A2(\wb_counter[5] ),
    .A3(_02336_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07544_ (.A1(\wb_counter[6] ),
    .A2(_02346_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07545_ (.A1(net390),
    .A2(_02344_),
    .B(_02330_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07546_ (.A1(_02341_),
    .A2(_02347_),
    .B(_02348_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07547_ (.A1(\wb_counter[4] ),
    .A2(\wb_counter[5] ),
    .A3(\wb_counter[6] ),
    .A4(_02336_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07548_ (.A1(\wb_counter[7] ),
    .A2(_02349_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07549_ (.I(_02292_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07550_ (.A1(net101),
    .A2(_02344_),
    .B(_02351_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07551_ (.A1(_02341_),
    .A2(_02350_),
    .B(_02352_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07552_ (.I(\wb_counter[7] ),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07553_ (.A1(_02353_),
    .A2(_02349_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07554_ (.A1(\wb_counter[8] ),
    .A2(_02354_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07555_ (.A1(net394),
    .A2(_02344_),
    .B(_02351_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07556_ (.A1(_02341_),
    .A2(_02355_),
    .B(_02356_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07557_ (.I(_02319_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07558_ (.I(_02357_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07559_ (.A1(\wb_counter[8] ),
    .A2(_02354_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07560_ (.A1(\wb_counter[9] ),
    .A2(_02359_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07561_ (.I(_02322_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07562_ (.A1(net404),
    .A2(_02361_),
    .B(_02351_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07563_ (.A1(_02358_),
    .A2(_02360_),
    .B(_02362_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07564_ (.A1(\wb_counter[9] ),
    .A2(_02359_),
    .B(\wb_counter[10] ),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07565_ (.A1(\wb_counter[9] ),
    .A2(\wb_counter[10] ),
    .A3(_02359_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07566_ (.A1(_02363_),
    .A2(_02364_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07567_ (.A1(net373),
    .A2(_02361_),
    .B(_02351_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07568_ (.A1(_02358_),
    .A2(_02365_),
    .B(net374),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07569_ (.A1(\wb_counter[11] ),
    .A2(_02364_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07570_ (.I(_02292_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07571_ (.A1(net377),
    .A2(_02361_),
    .B(_02368_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07572_ (.A1(_02358_),
    .A2(_02367_),
    .B(net378),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07573_ (.A1(\wb_counter[11] ),
    .A2(_02364_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07574_ (.A1(\wb_counter[12] ),
    .A2(_02370_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07575_ (.A1(net388),
    .A2(_02361_),
    .B(_02368_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07576_ (.A1(_02358_),
    .A2(_02371_),
    .B(_02372_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07577_ (.I(_02357_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07578_ (.A1(\wb_counter[11] ),
    .A2(\wb_counter[12] ),
    .A3(_02364_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07579_ (.A1(\wb_counter[13] ),
    .A2(_02374_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07580_ (.I(_02322_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07581_ (.A1(net396),
    .A2(_02376_),
    .B(_02368_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07582_ (.A1(_02373_),
    .A2(_02375_),
    .B(_02377_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07583_ (.I(\wb_counter[13] ),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07584_ (.A1(_02378_),
    .A2(_02374_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07585_ (.A1(\wb_counter[14] ),
    .A2(_02379_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07586_ (.A1(net398),
    .A2(_02376_),
    .B(_02368_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07587_ (.A1(_02373_),
    .A2(_02380_),
    .B(_02381_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07588_ (.A1(\wb_counter[14] ),
    .A2(_02379_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07589_ (.A1(\wb_counter[15] ),
    .A2(_02382_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07590_ (.I(_02073_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07591_ (.I(_02384_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07592_ (.A1(net402),
    .A2(_02376_),
    .B(_02385_),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07593_ (.A1(_02373_),
    .A2(_02383_),
    .B(_02386_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07594_ (.A1(\wb_counter[14] ),
    .A2(\wb_counter[15] ),
    .A3(_02379_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07595_ (.A1(\wb_counter[16] ),
    .A2(_02387_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07596_ (.A1(net386),
    .A2(_02376_),
    .B(_02385_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07597_ (.A1(_02373_),
    .A2(_02388_),
    .B(_02389_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07598_ (.I(_02357_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07599_ (.I(\wb_counter[16] ),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07600_ (.A1(_02391_),
    .A2(_02387_),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07601_ (.A1(\wb_counter[17] ),
    .A2(_02392_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07602_ (.I(_02339_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07603_ (.A1(net381),
    .A2(_02394_),
    .B(_02385_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07604_ (.A1(_02390_),
    .A2(_02393_),
    .B(net382),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07605_ (.A1(\wb_counter[17] ),
    .A2(_02392_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07606_ (.A1(\wb_counter[18] ),
    .A2(_02396_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07607_ (.A1(net81),
    .A2(_02394_),
    .B(_02385_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07608_ (.A1(_02390_),
    .A2(_02397_),
    .B(_02398_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07609_ (.A1(\wb_counter[17] ),
    .A2(\wb_counter[18] ),
    .A3(_02392_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07610_ (.A1(\wb_counter[19] ),
    .A2(_02399_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07611_ (.I(_02384_),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07612_ (.A1(net82),
    .A2(_02394_),
    .B(_02401_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07613_ (.A1(_02390_),
    .A2(_02400_),
    .B(_02402_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07614_ (.I(\wb_counter[19] ),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07615_ (.A1(_02403_),
    .A2(_02399_),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07616_ (.A1(\wb_counter[20] ),
    .A2(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07617_ (.A1(net84),
    .A2(_02394_),
    .B(_02401_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07618_ (.A1(_02390_),
    .A2(_02405_),
    .B(_02406_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07619_ (.I(_02357_),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07620_ (.A1(\wb_counter[20] ),
    .A2(_02404_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07621_ (.A1(\wb_counter[21] ),
    .A2(_02408_),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07622_ (.I(_02339_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07623_ (.A1(net85),
    .A2(_02410_),
    .B(_02401_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07624_ (.A1(_02407_),
    .A2(_02409_),
    .B(_02411_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07625_ (.A1(\wb_counter[20] ),
    .A2(\wb_counter[21] ),
    .A3(_02404_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07626_ (.A1(\wb_counter[22] ),
    .A2(_02412_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07627_ (.A1(net86),
    .A2(_02410_),
    .B(_02401_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07628_ (.A1(_02407_),
    .A2(_02413_),
    .B(_02414_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07629_ (.I(\wb_counter[22] ),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07630_ (.A1(_02415_),
    .A2(_02412_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07631_ (.A1(\wb_counter[23] ),
    .A2(_02416_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07632_ (.I(_02384_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07633_ (.A1(net87),
    .A2(_02410_),
    .B(_02418_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07634_ (.A1(_02407_),
    .A2(_02417_),
    .B(_02419_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07635_ (.A1(\wb_counter[23] ),
    .A2(_02416_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07636_ (.A1(\wb_counter[24] ),
    .A2(_02420_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07637_ (.A1(net88),
    .A2(_02410_),
    .B(_02418_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07638_ (.A1(_02407_),
    .A2(_02421_),
    .B(_02422_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07639_ (.I(_02320_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07640_ (.A1(\wb_counter[23] ),
    .A2(\wb_counter[24] ),
    .A3(_02416_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07641_ (.A1(\wb_counter[25] ),
    .A2(_02424_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07642_ (.I(_02339_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07643_ (.A1(net89),
    .A2(_02426_),
    .B(_02418_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07644_ (.A1(_02423_),
    .A2(_02425_),
    .B(_02427_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07645_ (.I(\wb_counter[25] ),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07646_ (.A1(_02428_),
    .A2(_02424_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07647_ (.A1(\wb_counter[26] ),
    .A2(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07648_ (.A1(net90),
    .A2(_02426_),
    .B(_02418_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07649_ (.A1(_02423_),
    .A2(_02430_),
    .B(_02431_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07650_ (.A1(\wb_counter[26] ),
    .A2(_02429_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07651_ (.A1(\wb_counter[27] ),
    .A2(_02432_),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07652_ (.I(_02384_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07653_ (.A1(net91),
    .A2(_02426_),
    .B(_02434_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07654_ (.A1(_02423_),
    .A2(_02433_),
    .B(_02435_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07655_ (.A1(\wb_counter[26] ),
    .A2(\wb_counter[27] ),
    .A3(_02429_),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07656_ (.A1(\wb_counter[28] ),
    .A2(_02436_),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07657_ (.A1(net92),
    .A2(_02426_),
    .B(_02434_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07658_ (.A1(_02423_),
    .A2(_02437_),
    .B(_02438_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07659_ (.I(\wb_counter[28] ),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07660_ (.A1(_02439_),
    .A2(_02436_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07661_ (.A1(\wb_counter[29] ),
    .A2(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07662_ (.A1(net392),
    .A2(_02340_),
    .B(_02434_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07663_ (.A1(_02332_),
    .A2(_02441_),
    .B(_02442_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07664_ (.A1(\wb_counter[29] ),
    .A2(_02440_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07665_ (.A1(\wb_counter[30] ),
    .A2(_02443_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07666_ (.A1(net400),
    .A2(_02340_),
    .B(_02434_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07667_ (.A1(_02332_),
    .A2(_02444_),
    .B(_02445_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07668_ (.A1(\wb_counter[29] ),
    .A2(\wb_counter[30] ),
    .A3(_02440_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07669_ (.A1(\wb_counter[31] ),
    .A2(_02446_),
    .Z(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07670_ (.A1(net96),
    .A2(_02340_),
    .B(_02074_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07671_ (.A1(_02332_),
    .A2(_02447_),
    .B(_02448_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07672_ (.I(_01538_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07673_ (.A1(net221),
    .A2(_01638_),
    .B(_01611_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07674_ (.A1(_02449_),
    .A2(_02450_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07675_ (.I(_01241_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07676_ (.I(_01550_),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07677_ (.A1(net228),
    .A2(_02452_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07678_ (.A1(_01055_),
    .A2(_01552_),
    .B(_02451_),
    .C(_02453_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07679_ (.A1(net248),
    .A2(net238),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07680_ (.A1(net229),
    .A2(_01628_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07681_ (.A1(_02454_),
    .A2(_02455_),
    .B(_02004_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07682_ (.A1(net230),
    .A2(_02452_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07683_ (.A1(_01060_),
    .A2(_01552_),
    .B(_02451_),
    .C(_02456_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07684_ (.A1(net231),
    .A2(_01638_),
    .B(_01654_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07685_ (.A1(_02449_),
    .A2(_02457_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07686_ (.A1(net232),
    .A2(_02452_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07687_ (.A1(_01067_),
    .A2(_01552_),
    .B(_02451_),
    .C(_02458_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07688_ (.A1(net252),
    .A2(net238),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07689_ (.A1(net233),
    .A2(_01628_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07690_ (.A1(_02459_),
    .A2(_02460_),
    .B(_02004_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07691_ (.A1(net234),
    .A2(_01628_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07692_ (.A1(_01038_),
    .A2(_02452_),
    .B(_02451_),
    .C(_02461_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07693_ (.I(_01723_),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07694_ (.A1(_02462_),
    .A2(_01534_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07695_ (.I(_01101_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07696_ (.I(_01577_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07697_ (.I(_02465_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07698_ (.I(_01281_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07699_ (.A1(_02467_),
    .A2(_01198_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07700_ (.I(_02468_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07701_ (.A1(_01276_),
    .A2(_01193_),
    .A3(_01216_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07702_ (.A1(_02469_),
    .A2(_02470_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07703_ (.A1(_02466_),
    .A2(_02471_),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07704_ (.I(_02472_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07705_ (.I(_01130_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07706_ (.A1(_01429_),
    .A2(_01224_),
    .A3(_01213_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07707_ (.A1(_01576_),
    .A2(_02475_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07708_ (.A1(_02474_),
    .A2(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07709_ (.I(_02477_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07710_ (.A1(_02473_),
    .A2(_02478_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07711_ (.A1(_02464_),
    .A2(_02479_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07712_ (.A1(_01943_),
    .A2(_02480_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07713_ (.I(_01274_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07714_ (.I(_02482_),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07715_ (.I(_02472_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07716_ (.I(_02484_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07717_ (.A1(\as2650.stack[3][13] ),
    .A2(_01693_),
    .B1(_01969_),
    .B2(\as2650.stack[2][13] ),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07718_ (.A1(_01873_),
    .A2(_01886_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07719_ (.I(_02487_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07720_ (.I(_02488_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07721_ (.I(_02489_),
    .Z(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07722_ (.I(_02490_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07723_ (.I(_02491_),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07724_ (.I(_02492_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07725_ (.A1(_01873_),
    .A2(\as2650.debug_psu[1] ),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07726_ (.I(_02494_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07727_ (.I(_02495_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07728_ (.I(_02496_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07729_ (.I(_02497_),
    .Z(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07730_ (.I(_02498_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07731_ (.I(_02499_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07732_ (.A1(\as2650.debug_psu[2] ),
    .A2(_01686_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07733_ (.I(_02501_),
    .Z(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07734_ (.I(_02502_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07735_ (.I(_02503_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07736_ (.I(_02504_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07737_ (.I(_02505_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07738_ (.A1(\as2650.stack[0][13] ),
    .A2(_02493_),
    .B1(_02500_),
    .B2(\as2650.stack[1][13] ),
    .C(_02506_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07739_ (.I(_01689_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07740_ (.I(_02508_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07741_ (.I(_02509_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07742_ (.I(_01965_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07743_ (.I(_02511_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07744_ (.I(_02512_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07745_ (.A1(\as2650.stack[7][13] ),
    .A2(_02510_),
    .B1(_02513_),
    .B2(\as2650.stack[6][13] ),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07746_ (.A1(\as2650.debug_psu[0] ),
    .A2(\as2650.debug_psu[1] ),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07747_ (.A1(\as2650.debug_psu[2] ),
    .A2(_02515_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07748_ (.I(_02516_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07749_ (.I(_02517_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07750_ (.I(_02518_),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07751_ (.I(_02519_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07752_ (.I(_02520_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07753_ (.A1(\as2650.stack[4][13] ),
    .A2(_02493_),
    .B1(_02500_),
    .B2(\as2650.stack[5][13] ),
    .C(_02521_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07754_ (.A1(_02486_),
    .A2(_02507_),
    .B1(_02514_),
    .B2(_02522_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07755_ (.A1(\as2650.stack[11][13] ),
    .A2(_01693_),
    .B1(_01969_),
    .B2(\as2650.stack[10][13] ),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07756_ (.I(_02489_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07757_ (.I(_02525_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07758_ (.I(_02526_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07759_ (.I(_02496_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07760_ (.I(_02528_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07761_ (.I(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07762_ (.A1(\as2650.stack[8][13] ),
    .A2(_02527_),
    .B1(_02530_),
    .B2(\as2650.stack[9][13] ),
    .C(_02506_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07763_ (.I(_02490_),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07764_ (.I(_02532_),
    .Z(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07765_ (.I(_02533_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07766_ (.I(_02497_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07767_ (.I(_02535_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07768_ (.I(_02536_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07769_ (.A1(\as2650.stack[12][13] ),
    .A2(_02534_),
    .B1(_02537_),
    .B2(\as2650.stack[13][13] ),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07770_ (.I(_02509_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07771_ (.I(_01965_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07772_ (.I(_02540_),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07773_ (.I(_02541_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07774_ (.A1(\as2650.stack[15][13] ),
    .A2(_02539_),
    .B1(_02542_),
    .B2(\as2650.stack[14][13] ),
    .C(_02521_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07775_ (.A1(_02524_),
    .A2(_02531_),
    .B1(_02538_),
    .B2(_02543_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07776_ (.A1(_01681_),
    .A2(\as2650.debug_psu[3] ),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07777_ (.A1(_01687_),
    .A2(_02545_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07778_ (.A1(_01681_),
    .A2(_02515_),
    .B(\as2650.debug_psu[3] ),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07779_ (.A1(_02546_),
    .A2(_02547_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07780_ (.I(_02548_),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07781_ (.I(_02549_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07782_ (.I(_02550_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07783_ (.I(_02551_),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _07784_ (.I0(_02523_),
    .I1(_02544_),
    .S(_02552_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07785_ (.I(_01172_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07786_ (.I(_01433_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07787_ (.A1(_02474_),
    .A2(_02554_),
    .A3(_02555_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07788_ (.I(_02556_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _07789_ (.A1(net216),
    .A2(_02485_),
    .B1(_02478_),
    .B2(_02553_),
    .C1(_02557_),
    .C2(_01462_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07790_ (.I(_02466_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07791_ (.I(_01459_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07792_ (.A1(_02560_),
    .A2(_01513_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07793_ (.A1(_01263_),
    .A2(_01244_),
    .A3(_02561_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07794_ (.A1(_01528_),
    .A2(_01151_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07795_ (.I(_02563_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07796_ (.A1(_02467_),
    .A2(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07797_ (.A1(_01183_),
    .A2(_02565_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07798_ (.I(_02566_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07799_ (.I(_02567_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07800_ (.A1(_02559_),
    .A2(_02562_),
    .A3(_02568_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07801_ (.I(_02569_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07802_ (.A1(_02483_),
    .A2(_02558_),
    .B(_02570_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07803_ (.I(_01254_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07804_ (.I(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07805_ (.A1(net63),
    .A2(net139),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07806_ (.A1(net139),
    .A2(_01157_),
    .B(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07807_ (.I(_02575_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07808_ (.I(_02576_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07809_ (.I(_01188_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07810_ (.I(_02578_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07811_ (.I(_02579_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07812_ (.A1(_01277_),
    .A2(_01364_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07813_ (.A1(_01204_),
    .A2(_01163_),
    .A3(_02581_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07814_ (.I(_02582_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07815_ (.A1(_01424_),
    .A2(_01508_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07816_ (.A1(_01233_),
    .A2(_01513_),
    .A3(_02583_),
    .A4(_02584_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07817_ (.I(_02585_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07818_ (.I(_02586_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07819_ (.A1(_02580_),
    .A2(_02561_),
    .A3(_02587_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07820_ (.A1(_01315_),
    .A2(_02588_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07821_ (.I(_01429_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07822_ (.A1(_02590_),
    .A2(_02576_),
    .B(_02567_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07823_ (.A1(_01092_),
    .A2(_02577_),
    .B(_02589_),
    .C(_02591_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07824_ (.A1(_02573_),
    .A2(_02592_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07825_ (.A1(_02481_),
    .A2(_02571_),
    .B(_02593_),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07826_ (.A1(_02463_),
    .A2(_02594_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07827_ (.I(_01574_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07828_ (.I(_02595_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07829_ (.A1(_01100_),
    .A2(_01286_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07830_ (.I(_02597_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07831_ (.I(_02598_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07832_ (.I(_02599_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _07833_ (.A1(_00681_),
    .A2(_00685_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07834_ (.I(_02601_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07835_ (.I(_02602_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07836_ (.I(_02462_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07837_ (.A1(\as2650.insin[0] ),
    .A2(_02596_),
    .B1(_02600_),
    .B2(_02603_),
    .C(_02604_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07838_ (.A1(_02449_),
    .A2(_02605_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _07839_ (.A1(_00667_),
    .A2(_00677_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07840_ (.I(_02606_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07841_ (.I(_02607_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07842_ (.A1(\as2650.insin[1] ),
    .A2(_02596_),
    .B1(_02600_),
    .B2(_02608_),
    .C(_02604_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07843_ (.A1(_02449_),
    .A2(_02609_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07844_ (.I(_01002_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07845_ (.I(_02610_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07846_ (.I(_01102_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07847_ (.A1(_01110_),
    .A2(_01112_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07848_ (.I(_02613_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07849_ (.I(_02614_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07850_ (.I(_02615_),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07851_ (.I(_02616_),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07852_ (.A1(\as2650.insin[2] ),
    .A2(_02612_),
    .B1(_02617_),
    .B2(_01288_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07853_ (.A1(_02611_),
    .A2(_02618_),
    .B(_02004_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07854_ (.I(_01124_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07855_ (.I(_02619_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07856_ (.A1(\as2650.insin[3] ),
    .A2(_02612_),
    .B1(_02620_),
    .B2(_01288_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07857_ (.I(_02003_),
    .Z(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07858_ (.A1(_02611_),
    .A2(_02621_),
    .B(_02622_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07859_ (.I(_01534_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07860_ (.I(_02623_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07861_ (.I(_01178_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07862_ (.I(_02625_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07863_ (.I(_02626_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07864_ (.I(_02627_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07865_ (.A1(\as2650.insin[4] ),
    .A2(_02596_),
    .B1(_02628_),
    .B2(_02600_),
    .C(_02604_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07866_ (.A1(_02624_),
    .A2(_02629_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07867_ (.I(_02462_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07868_ (.A1(\as2650.insin[5] ),
    .A2(_02596_),
    .B1(_02577_),
    .B2(_02600_),
    .C(_02630_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07869_ (.A1(_02624_),
    .A2(_02631_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07870_ (.I(_01334_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07871_ (.A1(_01319_),
    .A2(_01325_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07872_ (.A1(_01264_),
    .A2(_02633_),
    .A3(_01472_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07873_ (.I(_02634_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07874_ (.I(_01506_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07875_ (.I(_02636_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07876_ (.I(_01326_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07877_ (.I(_01721_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07878_ (.I(_02602_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07879_ (.A1(_02639_),
    .A2(_02640_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07880_ (.I(_01435_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07881_ (.I(_02642_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07882_ (.I(_02643_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07883_ (.I(_00686_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07884_ (.A1(_01720_),
    .A2(_02645_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07885_ (.I(_02643_),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07886_ (.A1(_02639_),
    .A2(_02647_),
    .B(_02602_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07887_ (.A1(_02644_),
    .A2(_02646_),
    .B(_02648_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07888_ (.A1(_02638_),
    .A2(_02641_),
    .B1(_02649_),
    .B2(_01320_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07889_ (.A1(_02637_),
    .A2(_01708_),
    .A3(_02650_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07890_ (.A1(\as2650.indirect_target[0] ),
    .A2(_02635_),
    .B(_02651_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07891_ (.I(_01294_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07892_ (.I(_02653_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07893_ (.A1(_01332_),
    .A2(_01304_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07894_ (.I(_02655_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07895_ (.I(_02656_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07896_ (.I(_02645_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07897_ (.I(_02658_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07898_ (.I(_01333_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07899_ (.I(_02660_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07900_ (.A1(_02659_),
    .A2(_02661_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07901_ (.A1(\as2650.indirect_target[0] ),
    .A2(_02654_),
    .B1(_02657_),
    .B2(_02662_),
    .C(_02463_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07902_ (.A1(_02632_),
    .A2(_02652_),
    .B(_02663_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07903_ (.A1(_01170_),
    .A2(_01300_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07904_ (.I(_01576_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07905_ (.A1(_01304_),
    .A2(_01483_),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07906_ (.I(_02666_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07907_ (.A1(_01427_),
    .A2(_02664_),
    .A3(_02665_),
    .A4(_02667_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07908_ (.I(_01546_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07909_ (.I(_02669_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07910_ (.A1(\as2650.cpu_hidden_rom_enable ),
    .A2(_02670_),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07911_ (.A1(\as2650.wb_hidden_rom_enable ),
    .A2(_01538_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07912_ (.A1(_02668_),
    .A2(_02671_),
    .B(_02672_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07913_ (.I(_01086_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07914_ (.I(_02673_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07915_ (.I(_00678_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07916_ (.I(_02675_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07917_ (.I(_02676_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07918_ (.I(_01702_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07919_ (.A1(_01264_),
    .A2(_02633_),
    .A3(_01472_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07920_ (.I(_02679_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07921_ (.A1(_00678_),
    .A2(_01743_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07922_ (.A1(_02646_),
    .A2(_02681_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07923_ (.I(_02642_),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07924_ (.A1(_02643_),
    .A2(_02682_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07925_ (.A1(_02607_),
    .A2(_02683_),
    .B(_02684_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07926_ (.A1(_01326_),
    .A2(_02682_),
    .B1(_02685_),
    .B2(_01319_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07927_ (.A1(_02000_),
    .A2(_02686_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07928_ (.A1(\as2650.indirect_target[1] ),
    .A2(_02680_),
    .B1(_02687_),
    .B2(_01453_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07929_ (.A1(_01251_),
    .A2(_01333_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07930_ (.A1(_02677_),
    .A2(_02678_),
    .A3(_02656_),
    .B1(_02688_),
    .B2(_02689_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07931_ (.A1(\as2650.indirect_target[1] ),
    .A2(_02573_),
    .B(_02690_),
    .C(_02630_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07932_ (.I(\as2650.irqs_latch[6] ),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07933_ (.I(\as2650.irqs_latch[2] ),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07934_ (.A1(\as2650.irqs_latch[1] ),
    .A2(_02693_),
    .B(\as2650.irqs_latch[3] ),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07935_ (.I(\as2650.irqs_latch[5] ),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07936_ (.A1(\as2650.irqs_latch[4] ),
    .A2(_02694_),
    .B(_02695_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07937_ (.A1(_02692_),
    .A2(_02696_),
    .B(\as2650.irqs_latch[7] ),
    .C(_01450_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07938_ (.A1(_02674_),
    .A2(_02691_),
    .A3(_02697_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07939_ (.I(_01334_),
    .Z(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07940_ (.A1(_01719_),
    .A2(_02645_),
    .A3(_02681_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07941_ (.A1(_02606_),
    .A2(_01744_),
    .B(_02699_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07942_ (.A1(_02615_),
    .A2(_01765_),
    .A3(_02700_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07943_ (.I(_02642_),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07944_ (.A1(_02702_),
    .A2(_02701_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07945_ (.A1(_02616_),
    .A2(_02644_),
    .B(_02703_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07946_ (.I(_01319_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07947_ (.A1(_02638_),
    .A2(_02701_),
    .B1(_02704_),
    .B2(_02705_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07948_ (.A1(_02001_),
    .A2(_02706_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07949_ (.I(_01468_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07950_ (.A1(_00611_),
    .A2(_02635_),
    .B1(_02707_),
    .B2(_02708_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07951_ (.A1(_02698_),
    .A2(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07952_ (.A1(_01250_),
    .A2(_01244_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07953_ (.I(_02711_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07954_ (.I(_02712_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07955_ (.A1(_01110_),
    .A2(_01112_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07956_ (.I(_02714_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07957_ (.I(_02715_),
    .Z(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07958_ (.A1(_02716_),
    .A2(_02678_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07959_ (.I(_02462_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07960_ (.A1(\as2650.indirect_target[2] ),
    .A2(_01259_),
    .B1(_02713_),
    .B2(_02717_),
    .C(_02718_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07961_ (.A1(\as2650.irqs_latch[4] ),
    .A2(\as2650.irqs_latch[5] ),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07962_ (.A1(\as2650.irqs_latch[2] ),
    .A2(\as2650.irqs_latch[3] ),
    .B(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07963_ (.A1(_01450_),
    .A2(\as2650.irqs_latch[6] ),
    .A3(\as2650.irqs_latch[7] ),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07964_ (.A1(_02710_),
    .A2(_02719_),
    .B1(_02721_),
    .B2(_02722_),
    .C(_01526_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07965_ (.I(_01305_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07966_ (.I(_02634_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07967_ (.A1(_01122_),
    .A2(_01123_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07968_ (.I(_02725_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07969_ (.A1(_02614_),
    .A2(_01764_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07970_ (.A1(_02614_),
    .A2(_01764_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07971_ (.A1(_02727_),
    .A2(_02700_),
    .B(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07972_ (.A1(_02726_),
    .A2(_01791_),
    .A3(_02729_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07973_ (.I(_02726_),
    .Z(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07974_ (.A1(_02643_),
    .A2(_02730_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07975_ (.A1(_02731_),
    .A2(_02702_),
    .B(_02732_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07976_ (.A1(_01326_),
    .A2(_02730_),
    .B1(_02733_),
    .B2(_02705_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(_02000_),
    .A2(_02734_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07978_ (.I(_01468_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07979_ (.A1(\as2650.indirect_target[3] ),
    .A2(_02724_),
    .B1(_02735_),
    .B2(_02736_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07980_ (.A1(_01335_),
    .A2(_02737_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07981_ (.I(_02731_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07982_ (.I(_02660_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07983_ (.I(_02711_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07984_ (.A1(_02739_),
    .A2(_02740_),
    .A3(_02741_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07985_ (.A1(\as2650.indirect_target[3] ),
    .A2(_02723_),
    .B(_02738_),
    .C(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07986_ (.I(_01450_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07987_ (.I(_02673_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07988_ (.A1(_02720_),
    .A2(_02722_),
    .B1(_02743_),
    .B2(_02744_),
    .C(_02745_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07989_ (.I(\as2650.ivectors_base[0] ),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07990_ (.I(_02718_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07991_ (.I(_01453_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07992_ (.A1(_02725_),
    .A2(_01791_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07993_ (.A1(_02725_),
    .A2(_01791_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07994_ (.A1(_02749_),
    .A2(_02729_),
    .B(_02750_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07995_ (.A1(_02626_),
    .A2(_01815_),
    .A3(_02751_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07996_ (.A1(_02647_),
    .A2(_02752_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07997_ (.A1(_02627_),
    .A2(_02644_),
    .B(_02753_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07998_ (.A1(_02638_),
    .A2(_02752_),
    .B1(_02754_),
    .B2(_01320_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07999_ (.A1(_02748_),
    .A2(_02001_),
    .A3(_02755_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08000_ (.I(_02679_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08001_ (.A1(\as2650.indirect_target[4] ),
    .A2(_02757_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08002_ (.A1(_02756_),
    .A2(_02758_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08003_ (.A1(_02632_),
    .A2(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08004_ (.I(_02572_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08005_ (.I(_02712_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08006_ (.I(_01153_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08007_ (.A1(_02763_),
    .A2(_01176_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08008_ (.A1(net62),
    .A2(_02763_),
    .B(_02764_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08009_ (.I(_02765_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08010_ (.A1(_02766_),
    .A2(_02678_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08011_ (.A1(\as2650.indirect_target[4] ),
    .A2(_02761_),
    .B1(_02762_),
    .B2(_02767_),
    .C(_02630_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08012_ (.A1(_02746_),
    .A2(_02747_),
    .B1(_02760_),
    .B2(_02768_),
    .C(_02745_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08013_ (.I(_01160_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08014_ (.I(_02769_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08015_ (.A1(_02625_),
    .A2(_01815_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08016_ (.A1(_02625_),
    .A2(_01815_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08017_ (.A1(_02771_),
    .A2(_02751_),
    .B(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08018_ (.A1(_02770_),
    .A2(_01829_),
    .A3(_02773_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08019_ (.A1(_02683_),
    .A2(_02774_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08020_ (.A1(_02770_),
    .A2(_02647_),
    .B(_02775_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08021_ (.A1(_02638_),
    .A2(_02774_),
    .B1(_02776_),
    .B2(_02705_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08022_ (.A1(_02000_),
    .A2(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08023_ (.A1(\as2650.indirect_target[5] ),
    .A2(_02635_),
    .B1(_02778_),
    .B2(_02708_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08024_ (.A1(_02698_),
    .A2(_02779_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08025_ (.I(_02770_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08026_ (.A1(_02781_),
    .A2(_02661_),
    .A3(_02741_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08027_ (.A1(\as2650.indirect_target[5] ),
    .A2(_02654_),
    .B(_02780_),
    .C(_02782_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08028_ (.A1(\as2650.ivectors_base[1] ),
    .A2(_02610_),
    .B(_01548_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08029_ (.A1(_02611_),
    .A2(_02783_),
    .B(_02784_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08030_ (.A1(_01153_),
    .A2(_01145_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08031_ (.A1(net64),
    .A2(_02763_),
    .B(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08032_ (.I(_02786_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08033_ (.I(_02787_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08034_ (.I(_02788_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08035_ (.I(_02789_),
    .Z(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08036_ (.I(_02790_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08037_ (.A1(_02791_),
    .A2(_02661_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08038_ (.A1(_02633_),
    .A2(_02683_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08039_ (.I(_02793_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08040_ (.A1(_02786_),
    .A2(_01845_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08041_ (.A1(_02769_),
    .A2(_01829_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08042_ (.A1(_01160_),
    .A2(_01829_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08043_ (.A1(_02796_),
    .A2(_02773_),
    .B(_02797_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08044_ (.A1(_02795_),
    .A2(_02798_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08045_ (.I(_01147_),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08046_ (.I(_02800_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08047_ (.I(_02801_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08048_ (.I(_02802_),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08049_ (.A1(_02803_),
    .A2(_02705_),
    .A3(_02647_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08050_ (.A1(_02794_),
    .A2(_02799_),
    .B(_02804_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08051_ (.A1(_02736_),
    .A2(_01456_),
    .A3(_02805_),
    .B1(_02724_),
    .B2(\as2650.indirect_target[6] ),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08052_ (.A1(_02698_),
    .A2(_02806_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08053_ (.A1(\as2650.indirect_target[6] ),
    .A2(_02654_),
    .B1(_02657_),
    .B2(_02792_),
    .C(_02807_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08054_ (.I(_01547_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08055_ (.A1(\as2650.ivectors_base[2] ),
    .A2(_02610_),
    .B(_02809_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08056_ (.A1(_02611_),
    .A2(_02808_),
    .B(_02810_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08057_ (.A1(_01153_),
    .A2(_01136_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08058_ (.A1(net65),
    .A2(_02763_),
    .B(_02811_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08059_ (.I(_02812_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08060_ (.I(_02813_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08061_ (.A1(_02814_),
    .A2(_02661_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08062_ (.A1(_02787_),
    .A2(_01864_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08063_ (.A1(_02795_),
    .A2(_02798_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08064_ (.A1(_02801_),
    .A2(_01845_),
    .B(_02817_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08065_ (.A1(_02816_),
    .A2(_02818_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08066_ (.A1(_02793_),
    .A2(_02819_),
    .B(_02804_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08067_ (.A1(_02736_),
    .A2(_01456_),
    .A3(_02820_),
    .B1(_02724_),
    .B2(\as2650.indirect_target[7] ),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08068_ (.A1(_01335_),
    .A2(_02821_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08069_ (.A1(\as2650.indirect_target[7] ),
    .A2(_02654_),
    .B1(_02657_),
    .B2(_02815_),
    .C(_02822_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08070_ (.A1(\as2650.ivectors_base[3] ),
    .A2(_02610_),
    .B(_02809_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08071_ (.A1(_02744_),
    .A2(_02823_),
    .B(_02824_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08072_ (.A1(_01877_),
    .A2(_01862_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08073_ (.A1(_01147_),
    .A2(_02825_),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08074_ (.I(_02786_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08075_ (.A1(_02827_),
    .A2(_01864_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08076_ (.A1(_02800_),
    .A2(_01845_),
    .B1(_02817_),
    .B2(_02816_),
    .C(_02828_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08077_ (.A1(_02826_),
    .A2(_02829_),
    .Z(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08078_ (.A1(_02794_),
    .A2(_02830_),
    .B(_02804_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08079_ (.A1(_02708_),
    .A2(_01456_),
    .A3(_02831_),
    .B1(_02724_),
    .B2(\as2650.indirect_target[8] ),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08080_ (.A1(\as2650.instruction_args_latch[8] ),
    .A2(_01702_),
    .A3(_02656_),
    .B1(\as2650.indirect_target[8] ),
    .B2(_02653_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08081_ (.A1(_02698_),
    .A2(_02832_),
    .B(_02833_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08082_ (.A1(_02604_),
    .A2(_02834_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08083_ (.A1(\as2650.ivectors_base[4] ),
    .A2(_02744_),
    .B(_02670_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08084_ (.A1(_02835_),
    .A2(_02836_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08085_ (.I(_02689_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08086_ (.A1(_02827_),
    .A2(_01892_),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08087_ (.A1(_02800_),
    .A2(_02825_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08088_ (.A1(_02839_),
    .A2(_02829_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08089_ (.A1(_02802_),
    .A2(_02825_),
    .B(_02840_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08090_ (.A1(_02838_),
    .A2(_02841_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08091_ (.A1(_02644_),
    .A2(_02634_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08092_ (.A1(_01258_),
    .A2(_02843_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08093_ (.A1(\as2650.indirect_target[9] ),
    .A2(_02757_),
    .B1(_02842_),
    .B2(_02844_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08094_ (.I(\as2650.instruction_args_latch[9] ),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08095_ (.A1(_02846_),
    .A2(_02740_),
    .A3(_02741_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08096_ (.I(_01723_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08097_ (.A1(\as2650.indirect_target[9] ),
    .A2(_01255_),
    .B(_02848_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08098_ (.A1(_02837_),
    .A2(_02845_),
    .B(_02847_),
    .C(_02849_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08099_ (.A1(\as2650.ivectors_base[5] ),
    .A2(_02744_),
    .B(_02850_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08100_ (.A1(_02624_),
    .A2(_02851_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08101_ (.I(_01002_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08102_ (.A1(_02787_),
    .A2(_01907_),
    .Z(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(_02801_),
    .A2(_01892_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08104_ (.A1(_02839_),
    .A2(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08105_ (.I(_02826_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08106_ (.A1(_02856_),
    .A2(_02829_),
    .A3(_02838_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08107_ (.A1(_02855_),
    .A2(_02857_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08108_ (.A1(_02853_),
    .A2(_02858_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08109_ (.A1(\as2650.indirect_target[10] ),
    .A2(_02680_),
    .B1(_02844_),
    .B2(_02859_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08110_ (.I(\as2650.instruction_args_latch[10] ),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08111_ (.A1(_02861_),
    .A2(_02740_),
    .A3(_02741_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08112_ (.A1(\as2650.indirect_target[10] ),
    .A2(_01255_),
    .B(_02848_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08113_ (.A1(_02837_),
    .A2(_02860_),
    .B(_02862_),
    .C(_02863_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08114_ (.A1(\as2650.ivectors_base[6] ),
    .A2(_02852_),
    .B(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08115_ (.A1(_02624_),
    .A2(_02865_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08116_ (.I(_02623_),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08117_ (.A1(_02800_),
    .A2(_01919_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08118_ (.A1(_02788_),
    .A2(_01908_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08119_ (.A1(_02868_),
    .A2(_02858_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08120_ (.A1(_02789_),
    .A2(_01908_),
    .B(_02869_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08121_ (.A1(_02867_),
    .A2(_02870_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08122_ (.A1(\as2650.indirect_target[11] ),
    .A2(_02680_),
    .B1(_02844_),
    .B2(_02871_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08123_ (.A1(\as2650.instruction_args_latch[11] ),
    .A2(_02740_),
    .A3(_02712_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08124_ (.A1(\as2650.indirect_target[11] ),
    .A2(_01330_),
    .B(_02848_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08125_ (.A1(_02837_),
    .A2(_02872_),
    .B(_02873_),
    .C(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08126_ (.A1(\as2650.ivectors_base[7] ),
    .A2(_02852_),
    .B(_02875_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08127_ (.A1(_02866_),
    .A2(_02876_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08128_ (.A1(_02788_),
    .A2(_01920_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08129_ (.A1(_02853_),
    .A2(_02867_),
    .Z(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08130_ (.A1(_02857_),
    .A2(_02878_),
    .B(_02855_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08131_ (.I0(_02789_),
    .I1(_02877_),
    .S(_02879_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08132_ (.A1(_02789_),
    .A2(_01908_),
    .B(_02880_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08133_ (.A1(_01936_),
    .A2(_02881_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08134_ (.A1(\as2650.indirect_target[12] ),
    .A2(_02680_),
    .B1(_02844_),
    .B2(_02882_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08135_ (.A1(\as2650.instruction_args_latch[12] ),
    .A2(_02660_),
    .A3(_02712_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08136_ (.A1(\as2650.indirect_target[12] ),
    .A2(_01330_),
    .B(_02848_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08137_ (.A1(_02837_),
    .A2(_02883_),
    .B(_02884_),
    .C(_02885_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08138_ (.A1(\as2650.ivectors_base[8] ),
    .A2(_02852_),
    .B(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08139_ (.A1(_02866_),
    .A2(_02887_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08140_ (.I(\as2650.ivectors_base[9] ),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08141_ (.A1(\as2650.indirect_target[13] ),
    .A2(_02757_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08142_ (.A1(_02636_),
    .A2(_00958_),
    .A3(_01708_),
    .A4(_02794_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08143_ (.A1(_02889_),
    .A2(_02890_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08144_ (.A1(_02632_),
    .A2(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08145_ (.I(\as2650.instruction_args_latch[13] ),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08146_ (.I(_02893_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08147_ (.I(_02894_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08148_ (.A1(_02895_),
    .A2(_01440_),
    .B(_02660_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08149_ (.A1(_00634_),
    .A2(_01440_),
    .B(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08150_ (.A1(\as2650.indirect_target[13] ),
    .A2(_02761_),
    .B1(_02713_),
    .B2(_02897_),
    .C(_02718_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08151_ (.A1(_02888_),
    .A2(_02747_),
    .B1(_02892_),
    .B2(_02898_),
    .C(_02745_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08152_ (.I(\as2650.ivectors_base[10] ),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08153_ (.A1(\as2650.indirect_target[14] ),
    .A2(_02757_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08154_ (.A1(_01949_),
    .A2(_02748_),
    .A3(_02001_),
    .A4(_02794_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08155_ (.A1(_02900_),
    .A2(_02901_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08156_ (.A1(_02632_),
    .A2(_02902_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08157_ (.I(_02572_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08158_ (.I(_00652_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08159_ (.A1(_01949_),
    .A2(_01298_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08160_ (.A1(_02905_),
    .A2(_01298_),
    .B(_02678_),
    .C(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08161_ (.A1(\as2650.indirect_target[14] ),
    .A2(_02904_),
    .B1(_02713_),
    .B2(_02907_),
    .C(_02718_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08162_ (.A1(_02899_),
    .A2(_02747_),
    .B1(_02903_),
    .B2(_02908_),
    .C(_02745_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08163_ (.A1(_02689_),
    .A2(_02635_),
    .B(_02653_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08164_ (.A1(_01335_),
    .A2(_02843_),
    .B(_00644_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08165_ (.A1(\as2650.indirect_target[15] ),
    .A2(_02909_),
    .B1(_02910_),
    .B2(_02723_),
    .C(_02630_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08166_ (.A1(\as2650.ivectors_base[11] ),
    .A2(_02852_),
    .B(_01548_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08167_ (.A1(_02911_),
    .A2(_02912_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _08168_ (.I(\as2650.instruction_args_latch[13] ),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08169_ (.A1(_02913_),
    .A2(_00652_),
    .B(_01296_),
    .C(_01722_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08170_ (.A1(_02713_),
    .A2(_02914_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08171_ (.A1(_01998_),
    .A2(\as2650.indexed_cyc[0] ),
    .A3(_02915_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08172_ (.A1(_01249_),
    .A2(_01242_),
    .A3(_02914_),
    .Z(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08173_ (.A1(_01748_),
    .A2(_02914_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08174_ (.I(_01167_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08175_ (.I(_02564_),
    .Z(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08176_ (.A1(_01130_),
    .A2(_02919_),
    .A3(_01206_),
    .A4(_02920_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08177_ (.A1(_02918_),
    .A2(_02921_),
    .B(_02664_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08178_ (.A1(_02895_),
    .A2(_02917_),
    .A3(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08179_ (.A1(_01292_),
    .A2(_01305_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08180_ (.A1(_01241_),
    .A2(_02924_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08181_ (.A1(_02916_),
    .A2(_02923_),
    .B(_02925_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08182_ (.A1(_01998_),
    .A2(\as2650.indexed_cyc[1] ),
    .A3(_02915_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08183_ (.I(\as2650.instruction_args_latch[14] ),
    .Z(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08184_ (.A1(_02927_),
    .A2(_02917_),
    .A3(_02922_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08185_ (.A1(_02926_),
    .A2(_02928_),
    .B(_02925_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08186_ (.A1(_01269_),
    .A2(_01320_),
    .B(_01334_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08187_ (.A1(_01998_),
    .A2(_01722_),
    .B1(_02653_),
    .B2(_02929_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08188_ (.A1(_01293_),
    .A2(_01306_),
    .B(_02930_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08189_ (.A1(_02747_),
    .A2(_02931_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08190_ (.A1(_02866_),
    .A2(_02932_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08191_ (.I(_01001_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08192_ (.A1(_01249_),
    .A2(_01297_),
    .A3(_01302_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08193_ (.I(_01336_),
    .Z(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08194_ (.A1(_02935_),
    .A2(_01202_),
    .A3(_01222_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08195_ (.I(_01265_),
    .Z(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08196_ (.A1(_01261_),
    .A2(_01298_),
    .A3(_01324_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08197_ (.A1(_01316_),
    .A2(_02938_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08198_ (.A1(_02937_),
    .A2(_02939_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08199_ (.A1(_02933_),
    .A2(_02934_),
    .A3(_02936_),
    .A4(_02940_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08200_ (.I(_01525_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08201_ (.A1(_01749_),
    .A2(_01223_),
    .B1(_02941_),
    .B2(_01295_),
    .C(_02942_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08202_ (.A1(_01221_),
    .A2(_02597_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08203_ (.I(_02943_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08204_ (.A1(_01233_),
    .A2(_02944_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08205_ (.A1(net213),
    .A2(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08206_ (.A1(_02866_),
    .A2(_02946_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08207_ (.I(\as2650.warmup[1] ),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08208_ (.A1(\as2650.warmup[0] ),
    .A2(_02947_),
    .B(_01034_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08209_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08210_ (.A1(_01034_),
    .A2(_02948_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08211_ (.I(_02623_),
    .Z(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08212_ (.I(_01485_),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08213_ (.A1(_01332_),
    .A2(_01308_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08214_ (.I(_02951_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08215_ (.A1(_01252_),
    .A2(_02603_),
    .B1(net195),
    .B2(_02952_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08216_ (.A1(_01336_),
    .A2(_01332_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08217_ (.I(_02954_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08218_ (.A1(_01040_),
    .A2(_02955_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08219_ (.A1(_02904_),
    .A2(_02953_),
    .B(_02956_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08220_ (.I(_02933_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08221_ (.A1(_01040_),
    .A2(_02950_),
    .B1(_02957_),
    .B2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08222_ (.A1(_02949_),
    .A2(_02959_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08223_ (.A1(_01252_),
    .A2(_02608_),
    .B1(net196),
    .B2(_02952_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08224_ (.A1(\as2650.instruction_args_latch[1] ),
    .A2(_02955_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08225_ (.A1(_02904_),
    .A2(_02960_),
    .B(_02961_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08226_ (.A1(\as2650.instruction_args_latch[1] ),
    .A2(_02950_),
    .B1(_02962_),
    .B2(_02958_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08227_ (.A1(_02949_),
    .A2(_02963_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08228_ (.A1(_01252_),
    .A2(_02617_),
    .B1(_02952_),
    .B2(net197),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08229_ (.A1(\as2650.instruction_args_latch[2] ),
    .A2(_02955_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08230_ (.A1(_02904_),
    .A2(_02964_),
    .B(_02965_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08231_ (.A1(\as2650.instruction_args_latch[2] ),
    .A2(_02950_),
    .B1(_02966_),
    .B2(_02958_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08232_ (.A1(_02949_),
    .A2(_02967_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08233_ (.I(_02572_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08234_ (.I(_01251_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08235_ (.A1(_02969_),
    .A2(_02620_),
    .B1(_02952_),
    .B2(net198),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08236_ (.A1(\as2650.instruction_args_latch[3] ),
    .A2(_02955_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08237_ (.A1(_02968_),
    .A2(_02970_),
    .B(_02971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08238_ (.A1(\as2650.instruction_args_latch[3] ),
    .A2(_02950_),
    .B1(_02972_),
    .B2(_02958_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08239_ (.A1(_02949_),
    .A2(_02973_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08240_ (.I(_02623_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08241_ (.I(_01485_),
    .Z(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08242_ (.I(_02951_),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08243_ (.A1(_02969_),
    .A2(_02628_),
    .B1(_02976_),
    .B2(net200),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08244_ (.I(_02954_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08245_ (.A1(\as2650.instruction_args_latch[4] ),
    .A2(_02978_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08246_ (.A1(_02968_),
    .A2(_02977_),
    .B(_02979_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08247_ (.I(_01001_),
    .Z(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08248_ (.A1(\as2650.instruction_args_latch[4] ),
    .A2(_02975_),
    .B1(_02980_),
    .B2(_02981_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08249_ (.A1(_02974_),
    .A2(_02982_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08250_ (.A1(_02969_),
    .A2(_02577_),
    .B1(_02976_),
    .B2(net201),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08251_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_02978_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08252_ (.A1(_02968_),
    .A2(_02983_),
    .B(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08253_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_02975_),
    .B1(_02985_),
    .B2(_02981_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08254_ (.A1(_02974_),
    .A2(_02986_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08255_ (.A1(_02969_),
    .A2(_02803_),
    .B1(_02976_),
    .B2(net202),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08256_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_02978_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08257_ (.A1(_02968_),
    .A2(_02987_),
    .B(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08258_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_02975_),
    .B1(_02989_),
    .B2(_02981_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08259_ (.A1(_02974_),
    .A2(_02990_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08260_ (.I(_01138_),
    .Z(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08261_ (.I(_02991_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08262_ (.A1(_01251_),
    .A2(_02992_),
    .B1(_02976_),
    .B2(net203),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08263_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_02978_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08264_ (.A1(_01259_),
    .A2(_02993_),
    .B(_02994_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08265_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_02975_),
    .B1(_02995_),
    .B2(_02981_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08266_ (.A1(_02974_),
    .A2(_02996_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08267_ (.I(_02933_),
    .Z(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08268_ (.I(_01480_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08269_ (.I(\as2650.instruction_args_latch[8] ),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08270_ (.I(_01265_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08271_ (.A1(_01506_),
    .A2(_01308_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08272_ (.I(_03001_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08273_ (.A1(_03000_),
    .A2(_02603_),
    .B1(net204),
    .B2(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08274_ (.A1(_02998_),
    .A2(_02637_),
    .A3(_02999_),
    .B1(_01259_),
    .B2(_03003_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08275_ (.A1(_02997_),
    .A2(_03004_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08276_ (.I(_01307_),
    .Z(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08277_ (.I(_03006_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08278_ (.A1(_03007_),
    .A2(\as2650.instruction_args_latch[8] ),
    .A3(_01256_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08279_ (.A1(_03005_),
    .A2(_03008_),
    .B(_02622_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08280_ (.I(_02846_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08281_ (.I(_01258_),
    .Z(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08282_ (.A1(_03000_),
    .A2(_02608_),
    .B1(net205),
    .B2(_03002_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08283_ (.A1(_02998_),
    .A2(_02637_),
    .A3(_03009_),
    .B1(_03010_),
    .B2(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08284_ (.A1(_02997_),
    .A2(_03012_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08285_ (.A1(_03007_),
    .A2(_02846_),
    .A3(_01256_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08286_ (.A1(_03013_),
    .A2(_03014_),
    .B(_02622_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08287_ (.A1(_03000_),
    .A2(_02617_),
    .B1(_03002_),
    .B2(net206),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08288_ (.A1(_03006_),
    .A2(_01315_),
    .A3(_02861_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08289_ (.A1(_02761_),
    .A2(_03015_),
    .B(_03016_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08290_ (.A1(_02997_),
    .A2(_03017_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08291_ (.A1(_03007_),
    .A2(_02861_),
    .A3(_01256_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08292_ (.A1(_03018_),
    .A2(_03019_),
    .B(_02622_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08293_ (.I(\as2650.instruction_args_latch[11] ),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08294_ (.I(_01265_),
    .Z(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08295_ (.I(_03001_),
    .Z(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08296_ (.A1(_03021_),
    .A2(_02620_),
    .B1(_03022_),
    .B2(net207),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08297_ (.A1(_02998_),
    .A2(_02637_),
    .A3(_03020_),
    .B1(_03010_),
    .B2(_03023_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08298_ (.A1(_02997_),
    .A2(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08299_ (.I(_01449_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08300_ (.A1(_03007_),
    .A2(\as2650.instruction_args_latch[11] ),
    .A3(_03026_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08301_ (.I(_02003_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08302_ (.A1(_03025_),
    .A2(_03027_),
    .B(_03028_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08303_ (.I(_02933_),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08304_ (.I(\as2650.instruction_args_latch[12] ),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08305_ (.A1(_03021_),
    .A2(_02627_),
    .B1(_03022_),
    .B2(net208),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08306_ (.A1(_02998_),
    .A2(_02937_),
    .A3(_03030_),
    .B1(_03010_),
    .B2(_03031_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08307_ (.A1(_03029_),
    .A2(_03032_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08308_ (.I(_03006_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08309_ (.A1(_03034_),
    .A2(\as2650.instruction_args_latch[12] ),
    .A3(_03026_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08310_ (.A1(_03033_),
    .A2(_03035_),
    .B(_03028_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08311_ (.I(_02913_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08312_ (.A1(_03021_),
    .A2(_02577_),
    .B1(_03022_),
    .B2(net209),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08313_ (.A1(_02935_),
    .A2(_02937_),
    .A3(_03036_),
    .B1(_03010_),
    .B2(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08314_ (.A1(_03029_),
    .A2(_03038_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08315_ (.A1(_03034_),
    .A2(_02895_),
    .A3(_03026_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08316_ (.A1(_03039_),
    .A2(_03040_),
    .B(_03028_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08317_ (.A1(_03021_),
    .A2(_02803_),
    .B1(_03022_),
    .B2(net211),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08318_ (.A1(_02935_),
    .A2(_02937_),
    .A3(_02905_),
    .B1(_01449_),
    .B2(_03041_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08319_ (.A1(_03029_),
    .A2(_03042_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08320_ (.A1(_03034_),
    .A2(_02927_),
    .A3(_03026_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08321_ (.A1(_03043_),
    .A2(_03044_),
    .B(_03028_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08322_ (.A1(_03000_),
    .A2(_02992_),
    .B1(_03002_),
    .B2(net212),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08323_ (.A1(_03006_),
    .A2(_01315_),
    .A3(_01299_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08324_ (.A1(_02761_),
    .A2(_03045_),
    .B(_03046_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08325_ (.A1(_03029_),
    .A2(_03047_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08326_ (.I(_01330_),
    .Z(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08327_ (.A1(_03034_),
    .A2(_01299_),
    .A3(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08328_ (.I(_01087_),
    .Z(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08329_ (.A1(_03048_),
    .A2(_03050_),
    .B(_03051_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08330_ (.A1(_02683_),
    .A2(_01474_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08331_ (.I(_03052_),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08332_ (.A1(_02636_),
    .A2(_00958_),
    .A3(_03053_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08333_ (.A1(_02934_),
    .A2(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08334_ (.A1(_02723_),
    .A2(_03055_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08335_ (.A1(_01131_),
    .A2(_02554_),
    .A3(_02555_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08336_ (.I(_03057_),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08337_ (.I(_03058_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08338_ (.A1(_01101_),
    .A2(_03059_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08339_ (.I(_03060_),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08340_ (.A1(_00634_),
    .A2(_03060_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08341_ (.A1(_01452_),
    .A2(_01475_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08342_ (.I(_03063_),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08343_ (.I(_03064_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08344_ (.A1(_02553_),
    .A2(_03061_),
    .B(_03062_),
    .C(_03065_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08345_ (.I(_01439_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08346_ (.A1(net212),
    .A2(_02991_),
    .A3(_03067_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08347_ (.A1(net211),
    .A2(_01438_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08348_ (.A1(_02788_),
    .A2(_03069_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08349_ (.A1(net209),
    .A2(_02575_),
    .A3(_03067_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08350_ (.A1(net208),
    .A2(_01437_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08351_ (.A1(_02765_),
    .A2(_03072_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08352_ (.A1(net207),
    .A2(_02619_),
    .A3(_01439_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08353_ (.A1(net206),
    .A2(_01436_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08354_ (.A1(_02714_),
    .A2(_03075_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08355_ (.A1(_02606_),
    .A2(net205),
    .A3(_01438_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08356_ (.A1(net205),
    .A2(_01436_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08357_ (.A1(_02675_),
    .A2(_03078_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08358_ (.A1(_02601_),
    .A2(_00844_),
    .A3(_01437_),
    .A4(_03079_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08359_ (.A1(_02614_),
    .A2(_03075_),
    .Z(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08360_ (.A1(_03077_),
    .A2(_03080_),
    .B(_03081_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08361_ (.A1(net207),
    .A2(_01437_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08362_ (.A1(_02725_),
    .A2(_03083_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08363_ (.A1(_03076_),
    .A2(_03082_),
    .B(_03084_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08364_ (.A1(_02625_),
    .A2(_03072_),
    .Z(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08365_ (.A1(_03074_),
    .A2(_03085_),
    .B(_03086_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08366_ (.A1(net209),
    .A2(_01438_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08367_ (.A1(_01160_),
    .A2(_03088_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08368_ (.A1(_03073_),
    .A2(_03087_),
    .B(_03089_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08369_ (.A1(_01147_),
    .A2(_03069_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08370_ (.A1(_03071_),
    .A2(_03090_),
    .B(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08371_ (.A1(net212),
    .A2(_01439_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08372_ (.A1(_02812_),
    .A2(_03093_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08373_ (.A1(_03070_),
    .A2(_03092_),
    .B(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08374_ (.A1(_03068_),
    .A2(_03095_),
    .B(_02999_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08375_ (.A1(\as2650.instruction_args_latch[9] ),
    .A2(\as2650.instruction_args_latch[10] ),
    .A3(_03096_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08376_ (.A1(_03020_),
    .A2(_03097_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08377_ (.A1(_03030_),
    .A2(_03098_),
    .Z(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08378_ (.A1(_02895_),
    .A2(_03099_),
    .Z(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08379_ (.A1(_01257_),
    .A2(_02934_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08380_ (.I(_03101_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08381_ (.I(_03102_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08382_ (.A1(_03056_),
    .A2(_03066_),
    .B1(_03100_),
    .B2(_03103_),
    .C(_02942_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08383_ (.I(_01240_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08384_ (.I(_03104_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08385_ (.A1(_01102_),
    .A2(_03059_),
    .B(_01949_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08386_ (.I(_02702_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08387_ (.I(_03063_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08388_ (.A1(\as2650.stack[3][14] ),
    .A2(_01693_),
    .B1(_01969_),
    .B2(\as2650.stack[2][14] ),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08389_ (.A1(\as2650.stack[0][14] ),
    .A2(_02493_),
    .B1(_02500_),
    .B2(\as2650.stack[1][14] ),
    .C(_02506_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08390_ (.A1(\as2650.stack[7][14] ),
    .A2(_02510_),
    .B1(_02513_),
    .B2(\as2650.stack[6][14] ),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08391_ (.A1(\as2650.stack[4][14] ),
    .A2(_02493_),
    .B1(_02500_),
    .B2(\as2650.stack[5][14] ),
    .C(_02521_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08392_ (.A1(_03109_),
    .A2(_03110_),
    .B1(_03111_),
    .B2(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08393_ (.A1(\as2650.stack[11][14] ),
    .A2(_02510_),
    .B1(_02513_),
    .B2(\as2650.stack[10][14] ),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08394_ (.A1(\as2650.stack[8][14] ),
    .A2(_02527_),
    .B1(_02530_),
    .B2(\as2650.stack[9][14] ),
    .C(_02506_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08395_ (.A1(\as2650.stack[12][14] ),
    .A2(_02534_),
    .B1(_02537_),
    .B2(\as2650.stack[13][14] ),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08396_ (.I(_02519_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08397_ (.A1(\as2650.stack[15][14] ),
    .A2(_02539_),
    .B1(_02542_),
    .B2(\as2650.stack[14][14] ),
    .C(_03117_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08398_ (.A1(_03114_),
    .A2(_03115_),
    .B1(_03116_),
    .B2(_03118_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08399_ (.I0(_03113_),
    .I1(_03119_),
    .S(_02552_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08400_ (.A1(_03107_),
    .A2(_03108_),
    .B1(_03120_),
    .B2(_03061_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08401_ (.A1(_03106_),
    .A2(_03121_),
    .B(_02667_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08402_ (.A1(_03036_),
    .A2(_02905_),
    .A3(_03099_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08403_ (.A1(_03036_),
    .A2(_03099_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08404_ (.A1(_02927_),
    .A2(_03124_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08405_ (.A1(_03123_),
    .A2(_03125_),
    .B(_03102_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08406_ (.A1(_03105_),
    .A2(_03122_),
    .A3(_03126_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08407_ (.I(_03127_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08408_ (.I(_02666_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08409_ (.A1(\as2650.stack[3][15] ),
    .A2(_02510_),
    .B1(_02513_),
    .B2(\as2650.stack[2][15] ),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08410_ (.I(_02503_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08411_ (.I(_03130_),
    .Z(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08412_ (.A1(\as2650.stack[0][15] ),
    .A2(_02527_),
    .B1(_02530_),
    .B2(\as2650.stack[1][15] ),
    .C(_03131_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08413_ (.A1(\as2650.stack[7][15] ),
    .A2(_02539_),
    .B1(_02542_),
    .B2(\as2650.stack[6][15] ),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08414_ (.A1(\as2650.stack[4][15] ),
    .A2(_02527_),
    .B1(_02530_),
    .B2(\as2650.stack[5][15] ),
    .C(_03117_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08415_ (.A1(_03129_),
    .A2(_03132_),
    .B1(_03133_),
    .B2(_03134_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08416_ (.A1(\as2650.stack[11][15] ),
    .A2(_02539_),
    .B1(_02542_),
    .B2(\as2650.stack[10][15] ),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08417_ (.I(_02532_),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08418_ (.I(_02535_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08419_ (.A1(\as2650.stack[8][15] ),
    .A2(_03137_),
    .B1(_03138_),
    .B2(\as2650.stack[9][15] ),
    .C(_03131_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08420_ (.A1(\as2650.stack[12][15] ),
    .A2(_02534_),
    .B1(_02537_),
    .B2(\as2650.stack[13][15] ),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08421_ (.I(_01691_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08422_ (.I(_01966_),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08423_ (.I(_03142_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08424_ (.A1(\as2650.stack[15][15] ),
    .A2(_03141_),
    .B1(_03143_),
    .B2(\as2650.stack[14][15] ),
    .C(_03117_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08425_ (.A1(_03136_),
    .A2(_03139_),
    .B1(_03140_),
    .B2(_03144_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08426_ (.I0(_03135_),
    .I1(_03145_),
    .S(_02552_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08427_ (.A1(_00644_),
    .A2(_03061_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08428_ (.A1(_03107_),
    .A2(_03065_),
    .B1(_03146_),
    .B2(_03061_),
    .C(_03147_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08429_ (.A1(_00649_),
    .A2(_03123_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08430_ (.A1(_03128_),
    .A2(_03149_),
    .B(_02809_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08431_ (.A1(_03128_),
    .A2(_03148_),
    .B(_03150_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08432_ (.A1(_01424_),
    .A2(_01282_),
    .A3(_01198_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08433_ (.A1(_03151_),
    .A2(_01578_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08434_ (.I(_02595_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08435_ (.A1(_02803_),
    .A2(_01337_),
    .B(_03152_),
    .C(_03153_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08436_ (.A1(\as2650.insin[6] ),
    .A2(_02612_),
    .B(_02463_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08437_ (.A1(_03154_),
    .A2(_03155_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08438_ (.A1(_02992_),
    .A2(_01337_),
    .B(_03152_),
    .C(_03153_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08439_ (.A1(\as2650.insin[7] ),
    .A2(_02612_),
    .B(_02463_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08440_ (.A1(_03156_),
    .A2(_03157_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08441_ (.I(_01727_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08442_ (.I(_01276_),
    .Z(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08443_ (.I(_01216_),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08444_ (.A1(_03158_),
    .A2(_03159_),
    .A3(_02579_),
    .A4(_03160_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08445_ (.A1(_02665_),
    .A2(_02943_),
    .A3(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08446_ (.I(_03162_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08447_ (.I(_03163_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08448_ (.I(_03163_),
    .Z(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08449_ (.A1(\as2650.ivectors_base[0] ),
    .A2(_03165_),
    .B(_02809_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08450_ (.A1(_01804_),
    .A2(_03164_),
    .B(_03166_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08451_ (.I(_01547_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08452_ (.A1(\as2650.ivectors_base[1] ),
    .A2(_03165_),
    .B(_03167_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08453_ (.A1(_01823_),
    .A2(_03164_),
    .B(_03168_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08454_ (.A1(\as2650.ivectors_base[2] ),
    .A2(_03165_),
    .B(_03167_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08455_ (.A1(_01838_),
    .A2(_03164_),
    .B(_03169_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08456_ (.A1(\as2650.ivectors_base[3] ),
    .A2(_03165_),
    .B(_03167_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08457_ (.A1(_01857_),
    .A2(_03164_),
    .B(_03170_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08458_ (.I(_03163_),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08459_ (.I(_03162_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08460_ (.A1(\as2650.ivectors_base[4] ),
    .A2(_03172_),
    .B(_03167_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08461_ (.A1(_01355_),
    .A2(_03171_),
    .B(_03173_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08462_ (.I(_01546_),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08463_ (.I(_03174_),
    .Z(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08464_ (.A1(\as2650.ivectors_base[5] ),
    .A2(_03172_),
    .B(_03175_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08465_ (.A1(_01351_),
    .A2(_03171_),
    .B(_03176_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08466_ (.A1(\as2650.ivectors_base[6] ),
    .A2(_03172_),
    .B(_03175_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08467_ (.A1(_01369_),
    .A2(_03171_),
    .B(_03177_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08468_ (.A1(\as2650.ivectors_base[7] ),
    .A2(_03172_),
    .B(_03175_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08469_ (.A1(_00831_),
    .A2(_03171_),
    .B(_03178_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08470_ (.I(_03163_),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08471_ (.I(_03162_),
    .Z(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08472_ (.A1(\as2650.ivectors_base[8] ),
    .A2(_03180_),
    .B(_03175_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08473_ (.A1(_00915_),
    .A2(_03179_),
    .B(_03181_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08474_ (.I(_03174_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08475_ (.A1(\as2650.ivectors_base[9] ),
    .A2(_03180_),
    .B(_03182_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08476_ (.A1(_00794_),
    .A2(_03179_),
    .B(_03183_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08477_ (.A1(\as2650.ivectors_base[10] ),
    .A2(_03180_),
    .B(_03182_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08478_ (.A1(_00774_),
    .A2(_03179_),
    .B(_03184_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08479_ (.A1(\as2650.ivectors_base[11] ),
    .A2(_03180_),
    .B(_03182_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08480_ (.A1(_00722_),
    .A2(_03179_),
    .B(_03185_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08481_ (.A1(_02640_),
    .A2(net204),
    .A3(_03067_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08482_ (.A1(net204),
    .A2(_03067_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08483_ (.A1(_02659_),
    .A2(_03187_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08484_ (.A1(_03186_),
    .A2(_03188_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08485_ (.I(_00597_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08486_ (.A1(_01297_),
    .A2(_01702_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08487_ (.I(_03191_),
    .Z(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08488_ (.A1(_03190_),
    .A2(_03192_),
    .B(_02655_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08489_ (.I(_03193_),
    .Z(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08490_ (.I(_03192_),
    .Z(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08491_ (.A1(_01721_),
    .A2(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08492_ (.I(_01274_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08493_ (.A1(_01219_),
    .A2(_01444_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08494_ (.A1(_03158_),
    .A2(_01217_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08495_ (.I(_01689_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08496_ (.A1(\as2650.stack[3][0] ),
    .A2(_03200_),
    .B1(_02511_),
    .B2(\as2650.stack[2][0] ),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08497_ (.A1(\as2650.stack[0][0] ),
    .A2(_02525_),
    .B1(_02528_),
    .B2(\as2650.stack[1][0] ),
    .C(_02504_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08498_ (.A1(\as2650.stack[7][0] ),
    .A2(_02508_),
    .B1(_02540_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08499_ (.I(_02517_),
    .Z(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08500_ (.A1(\as2650.stack[4][0] ),
    .A2(_02525_),
    .B1(_02528_),
    .B2(\as2650.stack[5][0] ),
    .C(_03204_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08501_ (.A1(_03201_),
    .A2(_03202_),
    .B1(_03203_),
    .B2(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08502_ (.A1(\as2650.stack[11][0] ),
    .A2(_03200_),
    .B1(_02511_),
    .B2(\as2650.stack[10][0] ),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08503_ (.A1(\as2650.stack[8][0] ),
    .A2(_02525_),
    .B1(_02528_),
    .B2(\as2650.stack[9][0] ),
    .C(_02504_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08504_ (.A1(\as2650.stack[12][0] ),
    .A2(_02532_),
    .B1(_02535_),
    .B2(\as2650.stack[13][0] ),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08505_ (.I(_01689_),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08506_ (.A1(\as2650.stack[15][0] ),
    .A2(_03210_),
    .B1(_02540_),
    .B2(\as2650.stack[14][0] ),
    .C(_03204_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08507_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03209_),
    .B2(_03211_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08508_ (.I0(_03206_),
    .I1(_03212_),
    .S(_02549_),
    .Z(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08509_ (.A1(_02554_),
    .A2(_02555_),
    .A3(_03213_),
    .B(_01219_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08510_ (.A1(_03198_),
    .A2(_03199_),
    .A3(_03214_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08511_ (.A1(_03197_),
    .A2(_03215_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08512_ (.A1(_02639_),
    .A2(_03216_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08513_ (.I(_03213_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08514_ (.A1(_02554_),
    .A2(_02555_),
    .A3(_03218_),
    .B(_01219_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08515_ (.A1(_03198_),
    .A2(_03199_),
    .A3(_03219_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08516_ (.A1(_01721_),
    .A2(_02482_),
    .A3(_03220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08517_ (.A1(_03217_),
    .A2(_03221_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08518_ (.A1(_00594_),
    .A2(_01473_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08519_ (.A1(_01452_),
    .A2(_03223_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08520_ (.I(_03224_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08521_ (.I(_01473_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08522_ (.A1(_01452_),
    .A2(_03226_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08523_ (.I(_03227_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08524_ (.I(_00641_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08525_ (.A1(_03229_),
    .A2(_02711_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08526_ (.A1(_02649_),
    .A2(_03064_),
    .B1(_03228_),
    .B2(_01045_),
    .C(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08527_ (.A1(_03222_),
    .A2(_03225_),
    .B(_03231_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08528_ (.A1(_03194_),
    .A2(_03196_),
    .B(_03232_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08529_ (.I(_02673_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08530_ (.A1(_03103_),
    .A2(_03189_),
    .B(_03233_),
    .C(_03234_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08531_ (.I(_03102_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08532_ (.A1(_03186_),
    .A2(_03079_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08533_ (.I(_03229_),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08534_ (.A1(_03237_),
    .A2(_01744_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08535_ (.A1(_03195_),
    .A2(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08536_ (.I(_03227_),
    .Z(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08537_ (.I(_03224_),
    .Z(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08538_ (.I(_01274_),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08539_ (.A1(_01443_),
    .A2(_03057_),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08540_ (.I(_03210_),
    .Z(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08541_ (.I(_01965_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08542_ (.I(_03245_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08543_ (.A1(\as2650.stack[3][1] ),
    .A2(_03244_),
    .B1(_03246_),
    .B2(\as2650.stack[2][1] ),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08544_ (.I(_02489_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08545_ (.I(_03248_),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08546_ (.I(_02496_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08547_ (.I(_03250_),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08548_ (.I(_02503_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08549_ (.A1(\as2650.stack[0][1] ),
    .A2(_03249_),
    .B1(_03251_),
    .B2(\as2650.stack[1][1] ),
    .C(_03252_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08550_ (.I(_03245_),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08551_ (.A1(\as2650.stack[7][1] ),
    .A2(_03244_),
    .B1(_03254_),
    .B2(\as2650.stack[6][1] ),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08552_ (.I(_02518_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08553_ (.A1(\as2650.stack[4][1] ),
    .A2(_03249_),
    .B1(_03251_),
    .B2(\as2650.stack[5][1] ),
    .C(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08554_ (.A1(_03247_),
    .A2(_03253_),
    .B1(_03255_),
    .B2(_03257_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08555_ (.A1(\as2650.stack[11][1] ),
    .A2(_03244_),
    .B1(_03246_),
    .B2(\as2650.stack[10][1] ),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08556_ (.A1(\as2650.stack[8][1] ),
    .A2(_03249_),
    .B1(_03251_),
    .B2(\as2650.stack[9][1] ),
    .C(_03252_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08557_ (.I(_03248_),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08558_ (.I(_03250_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08559_ (.A1(\as2650.stack[12][1] ),
    .A2(_03261_),
    .B1(_03262_),
    .B2(\as2650.stack[13][1] ),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08560_ (.I(_01690_),
    .Z(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08561_ (.A1(\as2650.stack[15][1] ),
    .A2(_03264_),
    .B1(_03254_),
    .B2(\as2650.stack[14][1] ),
    .C(_03256_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08562_ (.A1(_03259_),
    .A2(_03260_),
    .B1(_03263_),
    .B2(_03265_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08563_ (.I(_02549_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08564_ (.I0(_03258_),
    .I1(_03266_),
    .S(_03267_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08565_ (.A1(_01720_),
    .A2(_01128_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08566_ (.A1(_00606_),
    .A2(_03269_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08567_ (.A1(_01720_),
    .A2(_01762_),
    .A3(_01128_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08568_ (.A1(_01444_),
    .A2(_03270_),
    .A3(_03271_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08569_ (.A1(_01744_),
    .A2(_03243_),
    .B1(_03268_),
    .B2(_02557_),
    .C(_03272_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08570_ (.A1(_03242_),
    .A2(_03273_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08571_ (.A1(_01762_),
    .A2(_02482_),
    .B(_03241_),
    .C(_03274_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08572_ (.A1(_02685_),
    .A2(_03108_),
    .B1(_03240_),
    .B2(_03238_),
    .C(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08573_ (.I(_03230_),
    .Z(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08574_ (.I(_03277_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08575_ (.A1(_02762_),
    .A2(_03239_),
    .B1(_03276_),
    .B2(_03278_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08576_ (.A1(_03235_),
    .A2(_03236_),
    .B(_03279_),
    .C(_03234_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08577_ (.I(_03192_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08578_ (.A1(_03237_),
    .A2(_01765_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08579_ (.A1(_03280_),
    .A2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08580_ (.I(_01101_),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08581_ (.I(_01444_),
    .Z(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08582_ (.A1(_01789_),
    .A2(_03270_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08583_ (.A1(_00606_),
    .A2(_00610_),
    .A3(_03269_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08584_ (.A1(_03284_),
    .A2(_03285_),
    .A3(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08585_ (.A1(_01443_),
    .A2(_03057_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08586_ (.I(_01690_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08587_ (.I(_01966_),
    .Z(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08588_ (.A1(\as2650.stack[3][2] ),
    .A2(_03289_),
    .B1(_03290_),
    .B2(\as2650.stack[2][2] ),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08589_ (.I(_02490_),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08590_ (.I(_02497_),
    .Z(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08591_ (.I(_02503_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08592_ (.A1(\as2650.stack[0][2] ),
    .A2(_03292_),
    .B1(_03293_),
    .B2(\as2650.stack[1][2] ),
    .C(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08593_ (.I(_01966_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08594_ (.A1(\as2650.stack[7][2] ),
    .A2(_03289_),
    .B1(_03296_),
    .B2(\as2650.stack[6][2] ),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08595_ (.I(_02518_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08596_ (.A1(\as2650.stack[4][2] ),
    .A2(_03292_),
    .B1(_03293_),
    .B2(\as2650.stack[5][2] ),
    .C(_03298_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08597_ (.A1(_03291_),
    .A2(_03295_),
    .B1(_03297_),
    .B2(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08598_ (.A1(\as2650.stack[11][2] ),
    .A2(_03289_),
    .B1(_03290_),
    .B2(\as2650.stack[10][2] ),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08599_ (.I(_02490_),
    .Z(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08600_ (.I(_02497_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08601_ (.A1(\as2650.stack[8][2] ),
    .A2(_03302_),
    .B1(_03303_),
    .B2(\as2650.stack[9][2] ),
    .C(_03294_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08602_ (.I(_03248_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08603_ (.I(_03250_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08604_ (.A1(\as2650.stack[12][2] ),
    .A2(_03305_),
    .B1(_03306_),
    .B2(\as2650.stack[13][2] ),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08605_ (.I(_01690_),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08606_ (.A1(\as2650.stack[15][2] ),
    .A2(_03308_),
    .B1(_03142_),
    .B2(\as2650.stack[14][2] ),
    .C(_03298_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08607_ (.A1(_03301_),
    .A2(_03304_),
    .B1(_03307_),
    .B2(_03309_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08608_ (.I0(_03300_),
    .I1(_03310_),
    .S(_02550_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08609_ (.I(_03058_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08610_ (.A1(_01765_),
    .A2(_03288_),
    .B1(_03311_),
    .B2(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08611_ (.A1(_01275_),
    .A2(_03287_),
    .A3(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08612_ (.A1(_01789_),
    .A2(_03283_),
    .B(_03225_),
    .C(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08613_ (.A1(_02704_),
    .A2(_03108_),
    .B1(_03240_),
    .B2(_03281_),
    .C(_03315_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08614_ (.A1(_02762_),
    .A2(_03282_),
    .B1(_03316_),
    .B2(_03278_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08615_ (.A1(_03077_),
    .A2(_03080_),
    .A3(_03081_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08616_ (.A1(_03082_),
    .A2(_03318_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08617_ (.A1(_03128_),
    .A2(_03319_),
    .B(_01548_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08618_ (.A1(_03317_),
    .A2(_03320_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08619_ (.A1(_03076_),
    .A2(_03082_),
    .A3(_03084_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08620_ (.A1(_03085_),
    .A2(_03321_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08621_ (.A1(_01792_),
    .A2(_03195_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08622_ (.I(_03058_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08623_ (.A1(\as2650.stack[3][3] ),
    .A2(_03264_),
    .B1(_03254_),
    .B2(\as2650.stack[2][3] ),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08624_ (.A1(\as2650.stack[0][3] ),
    .A2(_03292_),
    .B1(_03293_),
    .B2(\as2650.stack[1][3] ),
    .C(_03252_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08625_ (.A1(\as2650.stack[7][3] ),
    .A2(_03264_),
    .B1(_03290_),
    .B2(\as2650.stack[6][3] ),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08626_ (.A1(\as2650.stack[4][3] ),
    .A2(_03305_),
    .B1(_03306_),
    .B2(\as2650.stack[5][3] ),
    .C(_03298_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08627_ (.A1(_03325_),
    .A2(_03326_),
    .B1(_03327_),
    .B2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08628_ (.A1(\as2650.stack[11][3] ),
    .A2(_03264_),
    .B1(_03290_),
    .B2(\as2650.stack[10][3] ),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08629_ (.A1(\as2650.stack[8][3] ),
    .A2(_03292_),
    .B1(_03293_),
    .B2(\as2650.stack[9][3] ),
    .C(_03294_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08630_ (.A1(\as2650.stack[12][3] ),
    .A2(_03305_),
    .B1(_03306_),
    .B2(\as2650.stack[13][3] ),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08631_ (.A1(\as2650.stack[15][3] ),
    .A2(_03308_),
    .B1(_03142_),
    .B2(\as2650.stack[14][3] ),
    .C(_03298_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08632_ (.A1(_03330_),
    .A2(_03331_),
    .B1(_03332_),
    .B2(_03333_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08633_ (.I0(_03329_),
    .I1(_03334_),
    .S(_03267_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08634_ (.A1(_00602_),
    .A2(_03285_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08635_ (.I(_01443_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08636_ (.A1(_03324_),
    .A2(_03335_),
    .B1(_03336_),
    .B2(_03337_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08637_ (.A1(_01792_),
    .A2(_03243_),
    .B(_03338_),
    .C(_03242_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08638_ (.A1(_01788_),
    .A2(_02464_),
    .B(_03339_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08639_ (.A1(_03229_),
    .A2(_01792_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08640_ (.A1(_02733_),
    .A2(_03064_),
    .B1(_03228_),
    .B2(_03341_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08641_ (.I(_03190_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08642_ (.A1(_03343_),
    .A2(_02655_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08643_ (.A1(_03225_),
    .A2(_03340_),
    .B(_03342_),
    .C(_03344_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08644_ (.A1(_03194_),
    .A2(_03323_),
    .B(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08645_ (.A1(_03235_),
    .A2(_03322_),
    .B(_03346_),
    .C(_03234_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08646_ (.I(_03191_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08647_ (.A1(_01816_),
    .A2(_03347_),
    .B(_03194_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08648_ (.A1(_01475_),
    .A2(_01816_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08649_ (.A1(_01475_),
    .A2(_02754_),
    .B1(_03349_),
    .B2(_03237_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08650_ (.I(_03288_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08651_ (.A1(\as2650.stack[3][4] ),
    .A2(_03289_),
    .B1(_03296_),
    .B2(\as2650.stack[2][4] ),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08652_ (.A1(\as2650.stack[0][4] ),
    .A2(_03302_),
    .B1(_03303_),
    .B2(\as2650.stack[1][4] ),
    .C(_03294_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08653_ (.A1(\as2650.stack[7][4] ),
    .A2(_03308_),
    .B1(_03296_),
    .B2(\as2650.stack[6][4] ),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08654_ (.A1(\as2650.stack[4][4] ),
    .A2(_03302_),
    .B1(_03303_),
    .B2(\as2650.stack[5][4] ),
    .C(_02519_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08655_ (.A1(_03352_),
    .A2(_03353_),
    .B1(_03354_),
    .B2(_03355_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08656_ (.A1(\as2650.stack[11][4] ),
    .A2(_03308_),
    .B1(_03296_),
    .B2(\as2650.stack[10][4] ),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08657_ (.A1(\as2650.stack[8][4] ),
    .A2(_03302_),
    .B1(_03303_),
    .B2(\as2650.stack[9][4] ),
    .C(_03130_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08658_ (.A1(\as2650.stack[12][4] ),
    .A2(_03305_),
    .B1(_03306_),
    .B2(\as2650.stack[13][4] ),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08659_ (.A1(\as2650.stack[15][4] ),
    .A2(_01691_),
    .B1(_01967_),
    .B2(\as2650.stack[14][4] ),
    .C(_02519_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08660_ (.A1(_03357_),
    .A2(_03358_),
    .B1(_03359_),
    .B2(_03360_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08661_ (.I0(_03356_),
    .I1(_03361_),
    .S(_02550_),
    .Z(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08662_ (.A1(_01789_),
    .A2(_01788_),
    .A3(_03270_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08663_ (.A1(_01813_),
    .A2(_03363_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08664_ (.A1(_03284_),
    .A2(_03364_),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08665_ (.A1(_01816_),
    .A2(_03351_),
    .B1(_03362_),
    .B2(_03059_),
    .C(_03365_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08666_ (.A1(_01812_),
    .A2(_01574_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08667_ (.A1(_02595_),
    .A2(_03366_),
    .B(_03367_),
    .C(_03225_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08668_ (.A1(_01469_),
    .A2(_03350_),
    .B(_03368_),
    .C(_03277_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08669_ (.A1(_03074_),
    .A2(_03085_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08670_ (.A1(_03086_),
    .A2(_03370_),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08671_ (.A1(_03348_),
    .A2(_03369_),
    .B1(_03371_),
    .B2(_03103_),
    .C(_02942_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08672_ (.I(_03193_),
    .Z(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08673_ (.A1(_01830_),
    .A2(_03280_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08674_ (.I(_03224_),
    .Z(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08675_ (.I(_03243_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08676_ (.A1(\as2650.stack[3][5] ),
    .A2(_01691_),
    .B1(_01967_),
    .B2(\as2650.stack[2][5] ),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08677_ (.A1(\as2650.stack[0][5] ),
    .A2(_02491_),
    .B1(_02498_),
    .B2(\as2650.stack[1][5] ),
    .C(_03130_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08678_ (.A1(\as2650.stack[7][5] ),
    .A2(_03200_),
    .B1(_02511_),
    .B2(\as2650.stack[6][5] ),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08679_ (.A1(\as2650.stack[4][5] ),
    .A2(_02491_),
    .B1(_02498_),
    .B2(\as2650.stack[5][5] ),
    .C(_03204_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08680_ (.A1(_03376_),
    .A2(_03377_),
    .B1(_03378_),
    .B2(_03379_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08681_ (.A1(\as2650.stack[11][5] ),
    .A2(_03200_),
    .B1(_01967_),
    .B2(\as2650.stack[10][5] ),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08682_ (.A1(\as2650.stack[8][5] ),
    .A2(_02491_),
    .B1(_02498_),
    .B2(\as2650.stack[9][5] ),
    .C(_03130_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08683_ (.A1(\as2650.stack[12][5] ),
    .A2(_02532_),
    .B1(_02535_),
    .B2(\as2650.stack[13][5] ),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08684_ (.A1(\as2650.stack[15][5] ),
    .A2(_02508_),
    .B1(_02540_),
    .B2(\as2650.stack[14][5] ),
    .C(_03204_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08685_ (.A1(_03381_),
    .A2(_03382_),
    .B1(_03383_),
    .B2(_03384_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08686_ (.I0(_03380_),
    .I1(_03385_),
    .S(_02550_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08687_ (.A1(_01813_),
    .A2(_03363_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08688_ (.A1(_01831_),
    .A2(_03387_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08689_ (.A1(_03324_),
    .A2(_03386_),
    .B1(_03388_),
    .B2(_01445_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08690_ (.A1(_01830_),
    .A2(_03375_),
    .B(_03389_),
    .C(_03197_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08691_ (.A1(_01831_),
    .A2(_03283_),
    .B(_03390_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08692_ (.A1(_03229_),
    .A2(_01830_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08693_ (.A1(_02776_),
    .A2(_03108_),
    .B1(_03228_),
    .B2(_03392_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08694_ (.A1(_03374_),
    .A2(_03391_),
    .B(_03393_),
    .C(_03344_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08695_ (.A1(_03372_),
    .A2(_03373_),
    .B(_03394_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08696_ (.A1(_03073_),
    .A2(_03087_),
    .A3(_03089_),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08697_ (.A1(_03090_),
    .A2(_03396_),
    .B(_02667_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08698_ (.A1(_02674_),
    .A2(_03395_),
    .A3(_03397_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08699_ (.A1(_01846_),
    .A2(_03347_),
    .B(_03372_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08700_ (.A1(_02802_),
    .A2(_02642_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08701_ (.A1(_03107_),
    .A2(_02799_),
    .B(_03399_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08702_ (.A1(_03343_),
    .A2(_01846_),
    .A3(_03240_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08703_ (.A1(_03344_),
    .A2(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08704_ (.I(_01574_),
    .Z(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08705_ (.A1(\as2650.stack[3][6] ),
    .A2(_01688_),
    .B1(_01964_),
    .B2(\as2650.stack[2][6] ),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08706_ (.A1(\as2650.stack[0][6] ),
    .A2(_02488_),
    .B1(_02495_),
    .B2(\as2650.stack[1][6] ),
    .C(_02502_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08707_ (.A1(\as2650.stack[7][6] ),
    .A2(_01688_),
    .B1(_01964_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08708_ (.A1(\as2650.stack[4][6] ),
    .A2(_02488_),
    .B1(_02495_),
    .B2(\as2650.stack[5][6] ),
    .C(_02516_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08709_ (.A1(_03404_),
    .A2(_03405_),
    .B1(_03406_),
    .B2(_03407_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08710_ (.A1(\as2650.stack[11][6] ),
    .A2(_01688_),
    .B1(_01964_),
    .B2(\as2650.stack[10][6] ),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08711_ (.A1(\as2650.stack[8][6] ),
    .A2(_02488_),
    .B1(_02495_),
    .B2(\as2650.stack[9][6] ),
    .C(_02501_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08712_ (.I(_02487_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08713_ (.I(_02494_),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08714_ (.A1(\as2650.stack[12][6] ),
    .A2(_03411_),
    .B1(_03412_),
    .B2(\as2650.stack[13][6] ),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08715_ (.A1(\as2650.stack[15][6] ),
    .A2(_01687_),
    .B1(_01963_),
    .B2(\as2650.stack[14][6] ),
    .C(_02516_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08716_ (.A1(_03409_),
    .A2(_03410_),
    .B1(_03413_),
    .B2(_03414_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08717_ (.I0(_03408_),
    .I1(_03415_),
    .S(_02548_),
    .Z(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08718_ (.A1(_01831_),
    .A2(_03387_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08719_ (.A1(_01848_),
    .A2(_03417_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08720_ (.A1(_03284_),
    .A2(_03418_),
    .Z(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08721_ (.A1(_01846_),
    .A2(_03351_),
    .B1(_03416_),
    .B2(_03059_),
    .C(_03419_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08722_ (.A1(_01848_),
    .A2(_02595_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08723_ (.A1(_03403_),
    .A2(_03420_),
    .B(_03421_),
    .C(_03374_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08724_ (.A1(_03065_),
    .A2(_03400_),
    .B(_03402_),
    .C(_03422_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08725_ (.A1(_03091_),
    .A2(_03071_),
    .A3(_03090_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08726_ (.A1(_03092_),
    .A2(_03424_),
    .B(_03101_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08727_ (.A1(_02670_),
    .A2(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08728_ (.A1(_03398_),
    .A2(_03423_),
    .B(_03426_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08729_ (.A1(_01865_),
    .A2(_03280_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08730_ (.I(_01687_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08731_ (.I(_01963_),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08732_ (.A1(\as2650.stack[3][7] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\as2650.stack[2][7] ),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08733_ (.A1(\as2650.stack[0][7] ),
    .A2(_03411_),
    .B1(_03412_),
    .B2(\as2650.stack[1][7] ),
    .C(_02502_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08734_ (.A1(\as2650.stack[7][7] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\as2650.stack[6][7] ),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08735_ (.A1(\as2650.stack[4][7] ),
    .A2(_03411_),
    .B1(_03412_),
    .B2(\as2650.stack[5][7] ),
    .C(_02517_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08736_ (.A1(_03430_),
    .A2(_03431_),
    .B1(_03432_),
    .B2(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08737_ (.A1(\as2650.stack[11][7] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\as2650.stack[10][7] ),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08738_ (.A1(\as2650.stack[8][7] ),
    .A2(_03411_),
    .B1(_03412_),
    .B2(\as2650.stack[9][7] ),
    .C(_02502_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08739_ (.A1(\as2650.stack[12][7] ),
    .A2(_02489_),
    .B1(_02496_),
    .B2(\as2650.stack[13][7] ),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08740_ (.A1(\as2650.stack[15][7] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\as2650.stack[14][7] ),
    .C(_02517_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08741_ (.A1(_03435_),
    .A2(_03436_),
    .B1(_03437_),
    .B2(_03438_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08742_ (.I0(_03434_),
    .I1(_03439_),
    .S(_02549_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08743_ (.A1(_01826_),
    .A2(_01848_),
    .A3(_03387_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08744_ (.A1(_00592_),
    .A2(_03441_),
    .Z(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08745_ (.A1(_03312_),
    .A2(_03440_),
    .B1(_03442_),
    .B2(_01445_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08746_ (.A1(_01865_),
    .A2(_03375_),
    .B(_03443_),
    .C(_03197_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08747_ (.A1(_01860_),
    .A2(_03283_),
    .B(_03444_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08748_ (.A1(_03237_),
    .A2(_01865_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08749_ (.A1(_03107_),
    .A2(_02819_),
    .B(_03399_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08750_ (.A1(_03228_),
    .A2(_03446_),
    .B1(_03447_),
    .B2(_03064_),
    .C(_03230_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08751_ (.A1(_03374_),
    .A2(_03445_),
    .B(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08752_ (.A1(_03372_),
    .A2(_03427_),
    .B(_03449_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08753_ (.A1(_03070_),
    .A2(_03092_),
    .A3(_03094_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08754_ (.A1(_03095_),
    .A2(_03451_),
    .B(_02667_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08755_ (.A1(_02674_),
    .A2(_03450_),
    .A3(_03452_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08756_ (.A1(_03068_),
    .A2(_03095_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08757_ (.A1(_02999_),
    .A2(_03453_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08758_ (.A1(_02702_),
    .A2(_02830_),
    .B(_03399_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08759_ (.A1(_00641_),
    .A2(_03226_),
    .A3(_01878_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08760_ (.A1(_03226_),
    .A2(_03455_),
    .B(_03456_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08761_ (.A1(_02825_),
    .A2(_03288_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08762_ (.A1(_00592_),
    .A2(_03441_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08763_ (.A1(_01879_),
    .A2(_03459_),
    .Z(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08764_ (.I(_03210_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08765_ (.I(_03245_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08766_ (.A1(\as2650.stack[3][8] ),
    .A2(_03461_),
    .B1(_03462_),
    .B2(\as2650.stack[2][8] ),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08767_ (.I(_02504_),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08768_ (.A1(\as2650.stack[0][8] ),
    .A2(_03261_),
    .B1(_03262_),
    .B2(\as2650.stack[1][8] ),
    .C(_03464_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08769_ (.I(_03210_),
    .Z(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08770_ (.A1(\as2650.stack[7][8] ),
    .A2(_03466_),
    .B1(_03462_),
    .B2(\as2650.stack[6][8] ),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08771_ (.A1(\as2650.stack[4][8] ),
    .A2(_03261_),
    .B1(_03262_),
    .B2(\as2650.stack[5][8] ),
    .C(_03256_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08772_ (.A1(_03463_),
    .A2(_03465_),
    .B1(_03467_),
    .B2(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08773_ (.A1(\as2650.stack[11][8] ),
    .A2(_03466_),
    .B1(_03462_),
    .B2(\as2650.stack[10][8] ),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08774_ (.A1(\as2650.stack[8][8] ),
    .A2(_03249_),
    .B1(_03251_),
    .B2(\as2650.stack[9][8] ),
    .C(_03252_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08775_ (.A1(\as2650.stack[12][8] ),
    .A2(_02526_),
    .B1(_02529_),
    .B2(\as2650.stack[13][8] ),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08776_ (.A1(\as2650.stack[15][8] ),
    .A2(_03244_),
    .B1(_03254_),
    .B2(\as2650.stack[14][8] ),
    .C(_03256_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08777_ (.A1(_03470_),
    .A2(_03471_),
    .B1(_03472_),
    .B2(_03473_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _08778_ (.I0(_03469_),
    .I1(_03474_),
    .S(_03267_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08779_ (.A1(_03337_),
    .A2(_03460_),
    .B1(_03475_),
    .B2(_03058_),
    .C(_01307_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08780_ (.A1(_01506_),
    .A2(_03457_),
    .B1(_03458_),
    .B2(_03476_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08781_ (.A1(_01879_),
    .A2(_02464_),
    .B1(_03477_),
    .B2(_01258_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08782_ (.A1(_03374_),
    .A2(_03457_),
    .B(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08783_ (.A1(_01878_),
    .A2(_03195_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08784_ (.A1(_03278_),
    .A2(_03479_),
    .B1(_03480_),
    .B2(_03194_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08785_ (.A1(_03235_),
    .A2(_03454_),
    .B(_03481_),
    .C(_03234_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08786_ (.A1(_01893_),
    .A2(_03347_),
    .B(_03193_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08787_ (.A1(_02636_),
    .A2(_03223_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08788_ (.A1(_01893_),
    .A2(_03351_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08789_ (.A1(_01879_),
    .A2(_03459_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08790_ (.A1(_01895_),
    .A2(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08791_ (.A1(\as2650.stack[3][9] ),
    .A2(_01692_),
    .B1(_02512_),
    .B2(\as2650.stack[2][9] ),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08792_ (.A1(\as2650.stack[0][9] ),
    .A2(_02492_),
    .B1(_02499_),
    .B2(\as2650.stack[1][9] ),
    .C(_02505_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08793_ (.A1(\as2650.stack[7][9] ),
    .A2(_02509_),
    .B1(_02512_),
    .B2(\as2650.stack[6][9] ),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08794_ (.A1(\as2650.stack[4][9] ),
    .A2(_02533_),
    .B1(_02536_),
    .B2(\as2650.stack[5][9] ),
    .C(_02520_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08795_ (.A1(_03487_),
    .A2(_03488_),
    .B1(_03489_),
    .B2(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08796_ (.A1(\as2650.stack[11][9] ),
    .A2(_02509_),
    .B1(_02512_),
    .B2(\as2650.stack[10][9] ),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08797_ (.A1(\as2650.stack[8][9] ),
    .A2(_02492_),
    .B1(_02499_),
    .B2(\as2650.stack[9][9] ),
    .C(_02505_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08798_ (.A1(\as2650.stack[12][9] ),
    .A2(_02533_),
    .B1(_02536_),
    .B2(\as2650.stack[13][9] ),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08799_ (.I(_02508_),
    .Z(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08800_ (.A1(\as2650.stack[15][9] ),
    .A2(_03495_),
    .B1(_02541_),
    .B2(\as2650.stack[14][9] ),
    .C(_02520_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08801_ (.A1(_03492_),
    .A2(_03493_),
    .B1(_03494_),
    .B2(_03496_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08802_ (.I0(_03491_),
    .I1(_03497_),
    .S(_02551_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08803_ (.A1(_01445_),
    .A2(_03486_),
    .B1(_03498_),
    .B2(_03312_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08804_ (.A1(_03197_),
    .A2(_03484_),
    .A3(_03499_),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08805_ (.A1(_01480_),
    .A2(_01895_),
    .B(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08806_ (.I(_03226_),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08807_ (.A1(_03502_),
    .A2(_01893_),
    .B1(_02842_),
    .B2(_03052_),
    .C(_03241_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08808_ (.A1(_03483_),
    .A2(_03501_),
    .B(_03503_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _08809_ (.A1(_01895_),
    .A2(_02723_),
    .B(_03277_),
    .C(_03504_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08810_ (.A1(_03009_),
    .A2(_03096_),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08811_ (.A1(_03482_),
    .A2(_03505_),
    .B1(_03506_),
    .B2(_03103_),
    .C(_02942_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08812_ (.A1(_02846_),
    .A2(_03096_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08813_ (.A1(_02861_),
    .A2(_03507_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08814_ (.A1(_03343_),
    .A2(_01909_),
    .B(_03192_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08815_ (.A1(_03190_),
    .A2(_01909_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08816_ (.A1(_02859_),
    .A2(_03053_),
    .B1(_03510_),
    .B2(_03502_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08817_ (.A1(_01877_),
    .A2(_01890_),
    .A3(_03459_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08818_ (.A1(_01917_),
    .A2(_03512_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08819_ (.I(_03245_),
    .Z(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08820_ (.A1(\as2650.stack[3][10] ),
    .A2(_03461_),
    .B1(_03514_),
    .B2(\as2650.stack[2][10] ),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08821_ (.I(_03248_),
    .Z(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08822_ (.I(_03250_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08823_ (.A1(\as2650.stack[0][10] ),
    .A2(_03516_),
    .B1(_03517_),
    .B2(\as2650.stack[1][10] ),
    .C(_03464_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08824_ (.A1(\as2650.stack[7][10] ),
    .A2(_03461_),
    .B1(_03462_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08825_ (.I(_02518_),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08826_ (.A1(\as2650.stack[4][10] ),
    .A2(_03516_),
    .B1(_03517_),
    .B2(\as2650.stack[5][10] ),
    .C(_03520_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08827_ (.A1(_03515_),
    .A2(_03518_),
    .B1(_03519_),
    .B2(_03521_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08828_ (.A1(\as2650.stack[11][10] ),
    .A2(_03461_),
    .B1(_03514_),
    .B2(\as2650.stack[10][10] ),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08829_ (.A1(\as2650.stack[8][10] ),
    .A2(_03261_),
    .B1(_03262_),
    .B2(\as2650.stack[9][10] ),
    .C(_03464_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08830_ (.A1(\as2650.stack[12][10] ),
    .A2(_02526_),
    .B1(_02529_),
    .B2(\as2650.stack[13][10] ),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08831_ (.A1(\as2650.stack[15][10] ),
    .A2(_03466_),
    .B1(_03246_),
    .B2(\as2650.stack[14][10] ),
    .C(_03520_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08832_ (.A1(_03523_),
    .A2(_03524_),
    .B1(_03525_),
    .B2(_03526_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08833_ (.I0(_03522_),
    .I1(_03527_),
    .S(_03267_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08834_ (.A1(_03337_),
    .A2(_03513_),
    .B1(_03528_),
    .B2(_03324_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08835_ (.A1(_01909_),
    .A2(_03375_),
    .B(_03529_),
    .C(_03242_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08836_ (.A1(_01905_),
    .A2(_02464_),
    .B(_03241_),
    .C(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08837_ (.A1(_01469_),
    .A2(_03511_),
    .B(_03531_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08838_ (.A1(_02762_),
    .A2(_03509_),
    .B1(_03532_),
    .B2(_03278_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08839_ (.I(_02673_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08840_ (.A1(_03235_),
    .A2(_03508_),
    .B(_03533_),
    .C(_03534_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08841_ (.A1(_01917_),
    .A2(_01916_),
    .A3(_03512_),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08842_ (.A1(_01917_),
    .A2(_03512_),
    .B(_01916_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08843_ (.A1(_03284_),
    .A2(_03535_),
    .A3(_03536_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08844_ (.A1(\as2650.stack[3][11] ),
    .A2(_03141_),
    .B1(_03143_),
    .B2(\as2650.stack[2][11] ),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08845_ (.A1(\as2650.stack[0][11] ),
    .A2(_03137_),
    .B1(_03138_),
    .B2(\as2650.stack[1][11] ),
    .C(_03131_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08846_ (.A1(\as2650.stack[7][11] ),
    .A2(_01692_),
    .B1(_01968_),
    .B2(\as2650.stack[6][11] ),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08847_ (.A1(\as2650.stack[4][11] ),
    .A2(_03137_),
    .B1(_03138_),
    .B2(\as2650.stack[5][11] ),
    .C(_03117_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08848_ (.A1(_03538_),
    .A2(_03539_),
    .B1(_03540_),
    .B2(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08849_ (.A1(\as2650.stack[11][11] ),
    .A2(_03141_),
    .B1(_01968_),
    .B2(\as2650.stack[10][11] ),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08850_ (.A1(\as2650.stack[8][11] ),
    .A2(_02533_),
    .B1(_02536_),
    .B2(\as2650.stack[9][11] ),
    .C(_03131_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08851_ (.A1(\as2650.stack[12][11] ),
    .A2(_03137_),
    .B1(_03138_),
    .B2(\as2650.stack[13][11] ),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08852_ (.A1(\as2650.stack[15][11] ),
    .A2(_01692_),
    .B1(_01968_),
    .B2(\as2650.stack[14][11] ),
    .C(_02520_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08853_ (.A1(_03543_),
    .A2(_03544_),
    .B1(_03545_),
    .B2(_03546_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08854_ (.I0(_03542_),
    .I1(_03547_),
    .S(_02551_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08855_ (.A1(_01920_),
    .A2(_03351_),
    .B1(_03548_),
    .B2(_03312_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08856_ (.A1(_01275_),
    .A2(_03537_),
    .A3(_03549_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08857_ (.A1(_02935_),
    .A2(_01915_),
    .B(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08858_ (.A1(_03190_),
    .A2(_01920_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08859_ (.A1(_02871_),
    .A2(_03053_),
    .B1(_03552_),
    .B2(_03502_),
    .C(_02736_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08860_ (.A1(_01916_),
    .A2(_01449_),
    .B1(_03483_),
    .B2(_03551_),
    .C(_03553_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08861_ (.A1(_03372_),
    .A2(_03554_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08862_ (.A1(_03098_),
    .A2(_03347_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08863_ (.A1(_03020_),
    .A2(_03097_),
    .B(_03556_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08864_ (.A1(_03280_),
    .A2(_03552_),
    .B(_03557_),
    .C(_02657_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08865_ (.A1(_02674_),
    .A2(_03555_),
    .A3(_03558_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08866_ (.A1(_03030_),
    .A2(_03098_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08867_ (.A1(_03099_),
    .A2(_03559_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08868_ (.A1(_02748_),
    .A2(_02882_),
    .A3(_03053_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08869_ (.A1(_01934_),
    .A2(_03535_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08870_ (.A1(\as2650.stack[3][12] ),
    .A2(_03495_),
    .B1(_02541_),
    .B2(\as2650.stack[2][12] ),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08871_ (.A1(\as2650.stack[0][12] ),
    .A2(_03516_),
    .B1(_03517_),
    .B2(\as2650.stack[1][12] ),
    .C(_02505_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08872_ (.A1(\as2650.stack[7][12] ),
    .A2(_03495_),
    .B1(_03514_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08873_ (.A1(\as2650.stack[4][12] ),
    .A2(_02526_),
    .B1(_02529_),
    .B2(\as2650.stack[5][12] ),
    .C(_03520_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08874_ (.A1(_03563_),
    .A2(_03564_),
    .B1(_03565_),
    .B2(_03566_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08875_ (.A1(\as2650.stack[11][12] ),
    .A2(_03495_),
    .B1(_02541_),
    .B2(\as2650.stack[10][12] ),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08876_ (.A1(\as2650.stack[8][12] ),
    .A2(_03516_),
    .B1(_03517_),
    .B2(\as2650.stack[9][12] ),
    .C(_03464_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08877_ (.A1(\as2650.stack[12][12] ),
    .A2(_02492_),
    .B1(_02499_),
    .B2(\as2650.stack[13][12] ),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08878_ (.A1(\as2650.stack[15][12] ),
    .A2(_03466_),
    .B1(_03246_),
    .B2(\as2650.stack[14][12] ),
    .C(_03520_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08879_ (.A1(_03568_),
    .A2(_03569_),
    .B1(_03570_),
    .B2(_03571_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08880_ (.I0(_03567_),
    .I1(_03572_),
    .S(_02551_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08881_ (.A1(_03337_),
    .A2(_03562_),
    .B1(_03573_),
    .B2(_03324_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08882_ (.A1(_01936_),
    .A2(_03375_),
    .B(_03574_),
    .C(_03242_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08883_ (.A1(_01934_),
    .A2(_03283_),
    .B(_03241_),
    .C(_03575_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08884_ (.A1(_03561_),
    .A2(_03576_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08885_ (.A1(_02656_),
    .A2(_03240_),
    .B(_03343_),
    .C(_01936_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08886_ (.A1(_03277_),
    .A2(_03577_),
    .B(_03578_),
    .C(_03101_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08887_ (.A1(_03102_),
    .A2(_03560_),
    .B(_03579_),
    .C(_03534_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08888_ (.I(\as2650.debug_psl[0] ),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08889_ (.A1(_01343_),
    .A2(_01227_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08890_ (.A1(_02812_),
    .A2(_01213_),
    .B(_03581_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08891_ (.A1(_01114_),
    .A2(_01209_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08892_ (.I(_03583_),
    .Z(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08893_ (.I(_03584_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08894_ (.I(_03585_),
    .Z(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08895_ (.I(_03586_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08896_ (.I(_03585_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08897_ (.I(_03588_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08898_ (.A1(_03589_),
    .A2(_01677_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08899_ (.A1(_01855_),
    .A2(_03587_),
    .B(_03590_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08900_ (.A1(_03582_),
    .A2(_03591_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08901_ (.A1(_01419_),
    .A2(_01212_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08902_ (.A1(_02786_),
    .A2(_01227_),
    .B(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08903_ (.A1(_03589_),
    .A2(_01669_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08904_ (.A1(_01667_),
    .A2(_03587_),
    .B(_03595_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08905_ (.A1(_03594_),
    .A2(_03596_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08906_ (.A1(_01346_),
    .A2(_01227_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08907_ (.A1(_02575_),
    .A2(_03589_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08908_ (.A1(_03598_),
    .A2(_03599_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08909_ (.A1(_03586_),
    .A2(_01660_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08910_ (.A1(_00803_),
    .A2(_03589_),
    .B(_03601_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08911_ (.A1(_03600_),
    .A2(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08912_ (.I(_03603_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08913_ (.A1(_01389_),
    .A2(_01211_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08914_ (.A1(_01178_),
    .A2(_03585_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _08915_ (.A1(_03605_),
    .A2(_03606_),
    .Z(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08916_ (.A1(_03588_),
    .A2(_01651_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08917_ (.A1(_00923_),
    .A2(_03586_),
    .B(_03608_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08918_ (.A1(_03607_),
    .A2(_03609_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08919_ (.A1(_00828_),
    .A2(_01226_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08920_ (.A1(_01124_),
    .A2(_03585_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08921_ (.A1(_03611_),
    .A2(_03612_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08922_ (.A1(_03588_),
    .A2(_01642_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08923_ (.A1(_00833_),
    .A2(_03586_),
    .B(_03614_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08924_ (.A1(_03613_),
    .A2(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08925_ (.A1(_01349_),
    .A2(_01225_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08926_ (.A1(_02613_),
    .A2(_03584_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08927_ (.A1(_03617_),
    .A2(_03618_),
    .Z(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08928_ (.A1(_01768_),
    .A2(_01211_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08929_ (.A1(_01211_),
    .A2(_01631_),
    .B(_03620_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08930_ (.A1(_03619_),
    .A2(_03621_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08931_ (.A1(_00881_),
    .A2(_01225_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08932_ (.A1(_02606_),
    .A2(_03583_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08933_ (.A1(_03623_),
    .A2(_03624_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08934_ (.I0(_01497_),
    .I1(_01620_),
    .S(_03584_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08935_ (.A1(_03625_),
    .A2(_03626_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08936_ (.A1(_01491_),
    .A2(_03584_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08937_ (.I(_01607_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08938_ (.A1(_00662_),
    .A2(_01373_),
    .B(_01225_),
    .C(_03629_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08939_ (.I0(_00686_),
    .I1(_01357_),
    .S(_01210_),
    .Z(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08940_ (.A1(_03628_),
    .A2(_03630_),
    .B(_03631_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08941_ (.A1(\as2650.debug_psl[0] ),
    .A2(\as2650.debug_psl[3] ),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08942_ (.I(_03633_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08943_ (.A1(_03631_),
    .A2(_03628_),
    .A3(_03630_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08944_ (.A1(_03632_),
    .A2(_03634_),
    .B(_03635_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08945_ (.A1(_03623_),
    .A2(_03624_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08946_ (.A1(_03637_),
    .A2(_03626_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08947_ (.A1(_03627_),
    .A2(_03636_),
    .B(_03638_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08948_ (.A1(_03611_),
    .A2(_03612_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08949_ (.A1(_00833_),
    .A2(_01226_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08950_ (.A1(_01212_),
    .A2(_01643_),
    .B(_03641_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08951_ (.A1(_03640_),
    .A2(_03642_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08952_ (.A1(_03619_),
    .A2(_03621_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08953_ (.A1(_03622_),
    .A2(_03639_),
    .B(_03643_),
    .C(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08954_ (.A1(_03605_),
    .A2(_03606_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08955_ (.I(_03609_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08956_ (.A1(_03646_),
    .A2(_03647_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08957_ (.A1(_03610_),
    .A2(_03616_),
    .A3(_03645_),
    .B(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08958_ (.I(_03602_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08959_ (.A1(_03600_),
    .A2(_03650_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08960_ (.A1(_03604_),
    .A2(_03649_),
    .B(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08961_ (.A1(_03594_),
    .A2(_03596_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08962_ (.A1(_03597_),
    .A2(_03652_),
    .B(_03653_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08963_ (.A1(_03582_),
    .A2(_03591_),
    .B(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08964_ (.A1(_01462_),
    .A2(_03592_),
    .A3(_03655_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08965_ (.I(_03582_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08966_ (.I(_00853_),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08967_ (.A1(_03658_),
    .A2(_01212_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _08968_ (.A1(_01606_),
    .A2(net356),
    .B(_03588_),
    .C(_01607_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08969_ (.I0(_02601_),
    .I1(_01373_),
    .S(_01226_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08970_ (.A1(_03659_),
    .A2(_03660_),
    .B(_03661_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08971_ (.A1(_01557_),
    .A2(_01779_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08972_ (.A1(_03635_),
    .A2(_03662_),
    .B(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08973_ (.A1(_03631_),
    .A2(_03659_),
    .A3(_03660_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08974_ (.I(_03626_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08975_ (.A1(_03637_),
    .A2(_03666_),
    .Z(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08976_ (.A1(_03664_),
    .A2(_03665_),
    .B(_03667_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08977_ (.A1(_03625_),
    .A2(_03666_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08978_ (.A1(_03617_),
    .A2(_03618_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08979_ (.I(_03621_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08980_ (.A1(_03670_),
    .A2(_03671_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08981_ (.A1(_03668_),
    .A2(_03669_),
    .B(_03672_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08982_ (.A1(_03670_),
    .A2(_03671_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08983_ (.I(_03616_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08984_ (.A1(_03675_),
    .A2(_03643_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08985_ (.A1(_03673_),
    .A2(_03674_),
    .B(_03676_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08986_ (.A1(_03613_),
    .A2(_03642_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08987_ (.I(_03610_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08988_ (.A1(_03677_),
    .A2(_03678_),
    .B(_03679_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08989_ (.A1(_03607_),
    .A2(_03647_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08990_ (.A1(_03600_),
    .A2(_03650_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08991_ (.A1(_03682_),
    .A2(_03604_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08992_ (.I(_03683_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08993_ (.A1(_03680_),
    .A2(_03681_),
    .B(_03684_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08994_ (.A1(_03598_),
    .A2(_03599_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08995_ (.A1(_03686_),
    .A2(_03650_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08996_ (.A1(_03594_),
    .A2(_03596_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08997_ (.A1(_03653_),
    .A2(_03688_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08998_ (.A1(_03685_),
    .A2(_03687_),
    .B(_03689_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _08999_ (.A1(_02787_),
    .A2(_01214_),
    .B(_03593_),
    .C(_03596_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09000_ (.I(_03592_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09001_ (.A1(_03582_),
    .A2(_03591_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09002_ (.A1(_03692_),
    .A2(_03693_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09003_ (.A1(_03690_),
    .A2(_03691_),
    .B(_03694_),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09004_ (.A1(_03657_),
    .A2(_03591_),
    .B(_03695_),
    .C(_01462_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09005_ (.A1(_02919_),
    .A2(_03696_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09006_ (.A1(_03580_),
    .A2(_02919_),
    .B1(_03656_),
    .B2(_03697_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09007_ (.I(_02587_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09008_ (.A1(_03699_),
    .A2(_02924_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09009_ (.A1(_01263_),
    .A2(_02561_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09010_ (.A1(_01257_),
    .A2(_03701_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09011_ (.I(_03702_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09012_ (.A1(_02466_),
    .A2(_02587_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09013_ (.I(_03704_),
    .Z(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09014_ (.I(_03580_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09015_ (.A1(_01183_),
    .A2(_02565_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09016_ (.I(_03707_),
    .Z(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09017_ (.I(_02590_),
    .Z(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09018_ (.A1(_03709_),
    .A2(_02602_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09019_ (.A1(_03706_),
    .A2(_02603_),
    .B(_03708_),
    .C(_03710_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09020_ (.A1(_03699_),
    .A2(_03698_),
    .B1(_03705_),
    .B2(_03711_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09021_ (.A1(_03703_),
    .A2(_03712_),
    .B(_03700_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09022_ (.A1(_01221_),
    .A2(_02598_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09023_ (.A1(_01232_),
    .A2(_01512_),
    .A3(_02582_),
    .A4(_02584_),
    .Z(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09024_ (.I(_03715_),
    .Z(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09025_ (.A1(_02579_),
    .A2(_02566_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09026_ (.I(_03717_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09027_ (.A1(_03716_),
    .A2(_03718_),
    .B(_03703_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09028_ (.I(_02578_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09029_ (.A1(_03720_),
    .A2(_02471_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09030_ (.I(_03721_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09031_ (.I(_03722_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09032_ (.A1(_01215_),
    .A2(_03716_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09033_ (.I(_03724_),
    .Z(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09034_ (.A1(_01195_),
    .A2(_02563_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09035_ (.A1(_01193_),
    .A2(_01215_),
    .A3(_03726_),
    .Z(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09036_ (.I(_03727_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09037_ (.I(_03587_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09038_ (.A1(_02474_),
    .A2(_03729_),
    .A3(_01367_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09039_ (.I(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09040_ (.I(_01779_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09041_ (.I(_03732_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09042_ (.A1(_03728_),
    .A2(_03731_),
    .B(_03733_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09043_ (.A1(_01575_),
    .A2(_02475_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09044_ (.A1(_01748_),
    .A2(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09045_ (.I(_03736_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09046_ (.A1(_03737_),
    .A2(_03218_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09047_ (.A1(_03706_),
    .A2(_03737_),
    .B(_03725_),
    .C(_03738_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09048_ (.A1(_03698_),
    .A2(_03725_),
    .B(_03734_),
    .C(_03739_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09049_ (.I(_01411_),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09050_ (.A1(_01193_),
    .A2(_01215_),
    .A3(_03726_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09051_ (.A1(_01204_),
    .A2(_01214_),
    .A3(_01398_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09052_ (.I(_01343_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09053_ (.I(_03744_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09054_ (.A1(_03741_),
    .A2(_03742_),
    .B1(_03743_),
    .B2(_03745_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09055_ (.I(_03721_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09056_ (.A1(_03733_),
    .A2(_03746_),
    .B(_03747_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09057_ (.A1(net188),
    .A2(_03723_),
    .B1(_03740_),
    .B2(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09058_ (.A1(_03714_),
    .A2(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09059_ (.A1(_03706_),
    .A2(_03714_),
    .B(_03719_),
    .C(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09060_ (.A1(_03698_),
    .A2(_03700_),
    .B1(_03713_),
    .B2(_03751_),
    .C(_01538_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09061_ (.I(_02003_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09062_ (.A1(_03703_),
    .A2(_03718_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09063_ (.I(_03737_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09064_ (.I(_03754_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09065_ (.A1(_03755_),
    .A2(_03268_),
    .B1(_03723_),
    .B2(net199),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09066_ (.A1(_03754_),
    .A2(_03747_),
    .B(_02482_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09067_ (.A1(_01755_),
    .A2(_03757_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09068_ (.A1(_03403_),
    .A2(_03756_),
    .B(_03758_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09069_ (.A1(_01755_),
    .A2(_02608_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09070_ (.A1(_00732_),
    .A2(_02677_),
    .B(_03708_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09071_ (.A1(_03701_),
    .A2(_03705_),
    .A3(_03760_),
    .A4(_03761_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09072_ (.A1(_03753_),
    .A2(_03759_),
    .B1(_03762_),
    .B2(_01295_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09073_ (.A1(_03752_),
    .A2(_03763_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09074_ (.A1(_02919_),
    .A2(_02586_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09075_ (.A1(_01293_),
    .A2(_03764_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09076_ (.A1(_03718_),
    .A2(_03764_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09077_ (.A1(_03701_),
    .A2(_03766_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09078_ (.A1(_01748_),
    .A2(_01703_),
    .A3(_02581_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09079_ (.I(_03768_),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09080_ (.A1(_03694_),
    .A2(_03690_),
    .A3(_03691_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09081_ (.A1(_03694_),
    .A2(_03654_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09082_ (.A1(_01698_),
    .A2(_01280_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09083_ (.I(_03772_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09084_ (.A1(_01197_),
    .A2(_01230_),
    .A3(_03772_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09085_ (.I(_03774_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09086_ (.I(_03775_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09087_ (.A1(_01283_),
    .A2(_03592_),
    .B(_03693_),
    .C(_02920_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09088_ (.A1(_03776_),
    .A2(_03777_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09089_ (.A1(_01169_),
    .A2(_03771_),
    .B1(_03773_),
    .B2(_03694_),
    .C(_03778_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09090_ (.A1(_01200_),
    .A2(_03695_),
    .A3(_03770_),
    .B(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09091_ (.A1(_03657_),
    .A2(_03776_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09092_ (.A1(_03780_),
    .A2(_03781_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09093_ (.I(_03782_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09094_ (.A1(_03592_),
    .A2(_03783_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09095_ (.A1(_03693_),
    .A2(_03783_),
    .B(_03784_),
    .C(_03764_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09096_ (.A1(_03729_),
    .A2(_02586_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09097_ (.A1(_03737_),
    .A2(_03311_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09098_ (.A1(_01771_),
    .A2(_02478_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09099_ (.A1(_01434_),
    .A2(_03786_),
    .B1(_03787_),
    .B2(_03788_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09100_ (.A1(_03722_),
    .A2(_03789_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09101_ (.A1(_03729_),
    .A2(_03769_),
    .A3(_03785_),
    .B(_03790_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09102_ (.A1(_01769_),
    .A2(_03747_),
    .B(_02944_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09103_ (.A1(_01772_),
    .A2(_02944_),
    .B1(_03791_),
    .B2(_03792_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09104_ (.A1(_03709_),
    .A2(_02615_),
    .B(_02567_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09105_ (.A1(_01771_),
    .A2(_02616_),
    .B(_03794_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09106_ (.A1(_03705_),
    .A2(_03795_),
    .B(_03785_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09107_ (.A1(_03702_),
    .A2(_03796_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09108_ (.A1(_03767_),
    .A2(_03793_),
    .B(_03797_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09109_ (.A1(_01292_),
    .A2(_01294_),
    .A3(_01513_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09110_ (.A1(_03769_),
    .A2(_03799_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09111_ (.I(_03785_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09112_ (.A1(_01772_),
    .A2(_03049_),
    .B1(_03765_),
    .B2(_03798_),
    .C1(_03800_),
    .C2(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09113_ (.A1(_03752_),
    .A2(_03802_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09114_ (.A1(_03755_),
    .A2(_03335_),
    .B1(_03723_),
    .B2(net214),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09115_ (.A1(_03733_),
    .A2(_03757_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09116_ (.A1(_03403_),
    .A2(_03803_),
    .B(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09117_ (.A1(_03753_),
    .A2(_03805_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09118_ (.A1(_03701_),
    .A2(_03705_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09119_ (.A1(_03159_),
    .A2(_02739_),
    .B(_03708_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09120_ (.A1(_01780_),
    .A2(_02739_),
    .B(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09121_ (.A1(_01295_),
    .A2(_03807_),
    .A3(_03809_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09122_ (.A1(_03806_),
    .A2(_03810_),
    .B(_03051_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09123_ (.A1(_03755_),
    .A2(_03362_),
    .B1(_03723_),
    .B2(net215),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09124_ (.I(_01807_),
    .Z(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09125_ (.I(_03812_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09126_ (.A1(_03813_),
    .A2(_03757_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09127_ (.A1(_03153_),
    .A2(_03811_),
    .B(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09128_ (.I(_01806_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09129_ (.I(_03816_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09130_ (.A1(_03709_),
    .A2(_02627_),
    .B(_02568_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09131_ (.A1(_03817_),
    .A2(_02628_),
    .B(_03807_),
    .C(_03818_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09132_ (.A1(_02573_),
    .A2(_03819_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09133_ (.A1(_03753_),
    .A2(_03815_),
    .B(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09134_ (.A1(_03752_),
    .A2(_03821_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09135_ (.A1(_01281_),
    .A2(_01166_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09136_ (.I(_03822_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09137_ (.I(_03610_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09138_ (.A1(_03661_),
    .A2(_03659_),
    .A3(_03660_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09139_ (.A1(\as2650.debug_psl[0] ),
    .A2(_01780_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09140_ (.A1(_03825_),
    .A2(_03632_),
    .B(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09141_ (.A1(_03661_),
    .A2(_03628_),
    .A3(_03630_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09142_ (.A1(_03827_),
    .A2(_03828_),
    .B(_03627_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09143_ (.A1(_03625_),
    .A2(_03666_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09144_ (.A1(_03829_),
    .A2(_03830_),
    .B(_03622_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09145_ (.A1(_03670_),
    .A2(_03671_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09146_ (.A1(_03616_),
    .A2(_03643_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09147_ (.A1(_03831_),
    .A2(_03832_),
    .B(_03833_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09148_ (.A1(_03640_),
    .A2(_03615_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09149_ (.A1(_03824_),
    .A2(_03834_),
    .A3(_03835_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09150_ (.A1(_03823_),
    .A2(_03680_),
    .A3(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09151_ (.A1(_03675_),
    .A2(_03645_),
    .B(_03679_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09152_ (.A1(_03679_),
    .A2(_03675_),
    .A3(_03645_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09153_ (.A1(_02469_),
    .A2(_03839_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09154_ (.A1(_01152_),
    .A2(_01195_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09155_ (.A1(_01167_),
    .A2(_02564_),
    .A3(_03841_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09156_ (.A1(_02467_),
    .A2(_03648_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09157_ (.A1(_03646_),
    .A2(_03647_),
    .B(_03843_),
    .C(_01231_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09158_ (.A1(_03679_),
    .A2(_03841_),
    .B(_03842_),
    .C(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09159_ (.A1(_03838_),
    .A2(_03840_),
    .B(_03845_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09160_ (.A1(_03607_),
    .A2(_03776_),
    .B1(_03837_),
    .B2(_03846_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09161_ (.A1(_03823_),
    .A2(_03824_),
    .A3(_03847_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09162_ (.A1(_03764_),
    .A2(_03848_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09163_ (.I(_03849_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09164_ (.A1(_01569_),
    .A2(_02478_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09165_ (.A1(_03736_),
    .A2(_03386_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09166_ (.A1(_01434_),
    .A2(_03786_),
    .B1(_03851_),
    .B2(_03852_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09167_ (.A1(_03160_),
    .A2(_03850_),
    .B(_03853_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09168_ (.I(_01419_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09169_ (.I(_03855_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09170_ (.I(_03856_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09171_ (.I(_01389_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09172_ (.A1(_03857_),
    .A2(_03742_),
    .B1(_03743_),
    .B2(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09173_ (.A1(_03734_),
    .A2(_03854_),
    .B1(_03859_),
    .B2(_03733_),
    .C(_03747_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09174_ (.A1(net216),
    .A2(_03722_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09175_ (.A1(_01336_),
    .A2(_01222_),
    .A3(_01337_),
    .A4(_03861_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09176_ (.A1(_01570_),
    .A2(_03714_),
    .B1(_03860_),
    .B2(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09177_ (.A1(_01569_),
    .A2(_02576_),
    .B(_02591_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09178_ (.A1(_03704_),
    .A2(_03864_),
    .B(_03849_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09179_ (.A1(_03702_),
    .A2(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09180_ (.A1(_03767_),
    .A2(_03863_),
    .B(_03866_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09181_ (.A1(_01570_),
    .A2(_03049_),
    .B1(_03800_),
    .B2(_03850_),
    .C1(_03867_),
    .C2(_03765_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09182_ (.A1(_03752_),
    .A2(_03868_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09183_ (.A1(_00765_),
    .A2(_00888_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09184_ (.A1(_01023_),
    .A2(_00816_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09185_ (.I(_00912_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09186_ (.A1(_01027_),
    .A2(_03871_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09187_ (.A1(_03872_),
    .A2(_03870_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09188_ (.A1(_03869_),
    .A2(_03873_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09189_ (.A1(_00790_),
    .A2(_00896_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09190_ (.A1(_00756_),
    .A2(_00874_),
    .B1(_00855_),
    .B2(_00717_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09191_ (.A1(_00717_),
    .A2(_00755_),
    .A3(_00874_),
    .A4(_00855_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09192_ (.A1(_03875_),
    .A2(_03876_),
    .B(_03877_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(_00754_),
    .A2(_00896_),
    .ZN(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09194_ (.A1(_00716_),
    .A2(_00873_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(_00790_),
    .A2(_00824_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09196_ (.A1(_03879_),
    .A2(_03880_),
    .A3(_03881_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09197_ (.A1(_03882_),
    .A2(_03878_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09198_ (.A1(_03878_),
    .A2(_03882_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09199_ (.A1(_03874_),
    .A2(_03883_),
    .B(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09200_ (.A1(_00728_),
    .A2(_00889_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09201_ (.A1(_00765_),
    .A2(_01013_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09202_ (.I(_01023_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09203_ (.A1(_03888_),
    .A2(_00914_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09204_ (.A1(_03886_),
    .A2(_03887_),
    .A3(_03889_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09205_ (.A1(_00757_),
    .A2(_01499_),
    .B1(_01494_),
    .B2(_00718_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09206_ (.I(_00755_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09207_ (.I(_01493_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09208_ (.A1(_00719_),
    .A2(_03892_),
    .A3(_01499_),
    .A4(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09209_ (.A1(_03881_),
    .A2(_03891_),
    .B(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09210_ (.A1(_00791_),
    .A2(_01028_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09211_ (.A1(_00755_),
    .A2(_00824_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09212_ (.A1(_00717_),
    .A2(_01498_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09213_ (.A1(_03896_),
    .A2(_03897_),
    .A3(_03898_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09214_ (.A1(_03895_),
    .A2(_03899_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09215_ (.A1(_03890_),
    .A2(_03900_),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09216_ (.A1(_03885_),
    .A2(_03901_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09217_ (.A1(_00767_),
    .A2(net189),
    .A3(_03873_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09218_ (.A1(_03870_),
    .A2(_03872_),
    .B(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09219_ (.A1(_03885_),
    .A2(_03901_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09220_ (.A1(_03904_),
    .A2(_03905_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09221_ (.I(_03886_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09222_ (.A1(_03887_),
    .A2(_03889_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09223_ (.A1(_03887_),
    .A2(_03889_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09224_ (.A1(_03907_),
    .A2(_03908_),
    .B(_03909_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09225_ (.A1(_03895_),
    .A2(_03899_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09226_ (.A1(_03890_),
    .A2(_03900_),
    .B(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09227_ (.A1(_00775_),
    .A2(_01012_),
    .B1(_01014_),
    .B2(_00729_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09228_ (.A1(_00728_),
    .A2(_00775_),
    .A3(_01012_),
    .A4(_01014_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09229_ (.I(_03914_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09230_ (.A1(_03913_),
    .A2(_03915_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09231_ (.A1(_03897_),
    .A2(_03898_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09232_ (.A1(_03897_),
    .A2(_03898_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09233_ (.A1(_03896_),
    .A2(_03917_),
    .B(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09234_ (.A1(_03892_),
    .A2(_01028_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09235_ (.A1(_00718_),
    .A2(_00826_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09236_ (.A1(_01023_),
    .A2(_00792_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09237_ (.A1(_03920_),
    .A2(_03921_),
    .A3(_03922_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09238_ (.A1(_03919_),
    .A2(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09239_ (.A1(_03916_),
    .A2(_03924_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09240_ (.A1(_03912_),
    .A2(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09241_ (.A1(_03910_),
    .A2(_03926_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09242_ (.A1(_03902_),
    .A2(_03906_),
    .B(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09243_ (.A1(_00728_),
    .A2(_01020_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09244_ (.A1(_01027_),
    .A2(_00888_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09245_ (.I(_00816_),
    .Z(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09246_ (.A1(_00826_),
    .A2(_03931_),
    .B1(_01498_),
    .B2(_00913_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09247_ (.A1(_00913_),
    .A2(_00825_),
    .A3(_03931_),
    .A4(_01498_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09248_ (.A1(_03930_),
    .A2(_03932_),
    .B(_03933_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09249_ (.A1(_00766_),
    .A2(_01016_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09250_ (.A1(_03934_),
    .A2(_03935_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09251_ (.A1(_03929_),
    .A2(_03936_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09252_ (.I(_00855_),
    .Z(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09253_ (.A1(_00756_),
    .A2(_00791_),
    .A3(_01493_),
    .A4(_03938_),
    .Z(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09254_ (.A1(_00824_),
    .A2(_00815_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09255_ (.A1(_03871_),
    .A2(_00897_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09256_ (.A1(_03930_),
    .A2(_03940_),
    .A3(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09257_ (.A1(_00792_),
    .A2(_00875_),
    .B1(_03938_),
    .B2(_03892_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09258_ (.A1(_03939_),
    .A2(_03942_),
    .A3(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09259_ (.A1(_00756_),
    .A2(_00791_),
    .A3(_01493_),
    .A4(_03938_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(_00754_),
    .A2(_00873_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09261_ (.A1(_00716_),
    .A2(_00854_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09262_ (.A1(_03946_),
    .A2(_03947_),
    .A3(_03875_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09263_ (.A1(_01022_),
    .A2(_00887_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09264_ (.A1(_01027_),
    .A2(_00815_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09265_ (.A1(_03871_),
    .A2(_00825_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09266_ (.A1(_03949_),
    .A2(_03950_),
    .A3(_03951_),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09267_ (.A1(_03945_),
    .A2(_03948_),
    .A3(_03952_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09268_ (.A1(_03953_),
    .A2(_03944_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09269_ (.A1(_03944_),
    .A2(_03953_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09270_ (.A1(_03937_),
    .A2(_03954_),
    .B(_03955_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09271_ (.A1(_03945_),
    .A2(_03948_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09272_ (.A1(_03945_),
    .A2(_03948_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09273_ (.A1(_03952_),
    .A2(_03957_),
    .B(_03958_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09274_ (.A1(_03874_),
    .A2(_03883_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09275_ (.A1(_03950_),
    .A2(_03951_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09276_ (.A1(_03950_),
    .A2(_03951_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09277_ (.A1(_03949_),
    .A2(_03961_),
    .B(_03962_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(_00729_),
    .A2(_01017_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09279_ (.A1(_03963_),
    .A2(_03964_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09280_ (.A1(_03959_),
    .A2(_03960_),
    .A3(_03965_),
    .Z(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09281_ (.A1(_03956_),
    .A2(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09282_ (.A1(net217),
    .A2(net220),
    .A3(_03934_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09283_ (.A1(_03929_),
    .A2(_03936_),
    .B(_03968_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09284_ (.A1(_03966_),
    .A2(_03956_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09285_ (.A1(_03969_),
    .A2(_03970_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09286_ (.A1(_03967_),
    .A2(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09287_ (.A1(_03963_),
    .A2(_03964_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09288_ (.I(_03965_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09289_ (.A1(_03959_),
    .A2(_03960_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09290_ (.A1(_03959_),
    .A2(_03960_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09291_ (.A1(_03974_),
    .A2(_03975_),
    .B(_03976_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09292_ (.A1(_03904_),
    .A2(_03905_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09293_ (.A1(_03978_),
    .A2(_03977_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09294_ (.A1(_03973_),
    .A2(_03979_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09295_ (.A1(_03972_),
    .A2(_03980_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(_00766_),
    .A2(_01019_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09297_ (.A1(_00825_),
    .A2(_00888_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09298_ (.A1(_01013_),
    .A2(_00898_),
    .B1(_00875_),
    .B2(_00913_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09299_ (.I(_03871_),
    .Z(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09300_ (.A1(_03985_),
    .A2(_03931_),
    .A3(_00898_),
    .A4(_00875_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09301_ (.A1(_03983_),
    .A2(_03984_),
    .B(_03986_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09302_ (.A1(_01024_),
    .A2(_01016_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09303_ (.A1(_03987_),
    .A2(_03988_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09304_ (.A1(_01024_),
    .A2(net220),
    .A3(_03987_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09305_ (.A1(_03982_),
    .A2(_03989_),
    .B(_03990_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09306_ (.A1(_03982_),
    .A2(_03989_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09307_ (.A1(_00792_),
    .A2(_00856_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09308_ (.A1(_03931_),
    .A2(_00897_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09309_ (.A1(_03985_),
    .A2(_03893_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09310_ (.A1(_03983_),
    .A2(_03994_),
    .A3(_03995_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09311_ (.A1(_03993_),
    .A2(_03996_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09312_ (.A1(_03939_),
    .A2(_03943_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09313_ (.A1(_03942_),
    .A2(_03998_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09314_ (.A1(_03997_),
    .A2(_03999_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(_03997_),
    .A2(_03999_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09316_ (.A1(_03992_),
    .A2(_04000_),
    .B(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09317_ (.A1(_03937_),
    .A2(_03954_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09318_ (.A1(_04002_),
    .A2(_04003_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09319_ (.A1(_04002_),
    .A2(_04003_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09320_ (.A1(_03991_),
    .A2(_04004_),
    .B(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09321_ (.A1(_03969_),
    .A2(_03970_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09322_ (.A1(_04006_),
    .A2(_04007_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09323_ (.A1(_01029_),
    .A2(_01019_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09324_ (.A1(_00826_),
    .A2(_01016_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09325_ (.A1(_01014_),
    .A2(_01015_),
    .A3(_01494_),
    .A4(_01489_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09326_ (.A1(_04009_),
    .A2(_04010_),
    .A3(_04011_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09327_ (.A1(_00817_),
    .A2(_01494_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(_00914_),
    .A2(_01489_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09329_ (.A1(_00898_),
    .A2(_00889_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09330_ (.A1(_04013_),
    .A2(_04014_),
    .A3(_04015_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09331_ (.A1(_04012_),
    .A2(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09332_ (.A1(_01499_),
    .A2(_01017_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09333_ (.A1(_01501_),
    .A2(_01020_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09334_ (.A1(_04018_),
    .A2(_04019_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09335_ (.A1(_01015_),
    .A2(_01495_),
    .B1(_01489_),
    .B2(net190),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09336_ (.A1(_04011_),
    .A2(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09337_ (.A1(_04018_),
    .A2(_04019_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09338_ (.A1(_04020_),
    .A2(_04022_),
    .B(_04023_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09339_ (.A1(_04017_),
    .A2(_04024_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09340_ (.A1(_01015_),
    .A2(_01490_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09341_ (.I(_01020_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09342_ (.A1(_01496_),
    .A2(_01018_),
    .B1(_04027_),
    .B2(_01500_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09343_ (.A1(_01500_),
    .A2(_01495_),
    .A3(_01018_),
    .A4(_04027_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09344_ (.A1(_04026_),
    .A2(_04028_),
    .B(_04029_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09345_ (.A1(_04020_),
    .A2(_04022_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09346_ (.A1(_04030_),
    .A2(_04031_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09347_ (.A1(_01500_),
    .A2(_04027_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09348_ (.A1(_01495_),
    .A2(_01018_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09349_ (.A1(_04033_),
    .A2(_04034_),
    .A3(_04026_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09350_ (.A1(_01496_),
    .A2(_04027_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09351_ (.A1(net220),
    .A2(_01490_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09352_ (.A1(_04036_),
    .A2(_04037_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09353_ (.A1(_04035_),
    .A2(_04038_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09354_ (.A1(_04020_),
    .A2(_04022_),
    .A3(_04030_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09355_ (.A1(_04039_),
    .A2(_04040_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09356_ (.A1(_04017_),
    .A2(_04024_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09357_ (.A1(_04032_),
    .A2(_04041_),
    .B(_04042_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09358_ (.A1(_04010_),
    .A2(_04011_),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09359_ (.A1(_01030_),
    .A2(_01021_),
    .A3(_04044_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09360_ (.A1(_04010_),
    .A2(_04011_),
    .B(_04045_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09361_ (.A1(_03993_),
    .A2(_03996_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09362_ (.A1(_03888_),
    .A2(_01019_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09363_ (.A1(_00817_),
    .A2(_03893_),
    .B1(_03938_),
    .B2(_03985_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09364_ (.A1(_03985_),
    .A2(_01013_),
    .A3(_03893_),
    .A4(_00856_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09365_ (.A1(_04015_),
    .A2(_04049_),
    .B(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09366_ (.A1(_01029_),
    .A2(_01017_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09367_ (.A1(_04048_),
    .A2(_04051_),
    .A3(_04052_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09368_ (.A1(_04012_),
    .A2(_04016_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09369_ (.A1(_04047_),
    .A2(_04053_),
    .A3(_04054_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09370_ (.A1(_04046_),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09371_ (.A1(_04025_),
    .A2(_04043_),
    .B(_04056_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09372_ (.A1(_04047_),
    .A2(_04053_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09373_ (.A1(_04012_),
    .A2(_04016_),
    .A3(_04058_),
    .B1(_04046_),
    .B2(_04055_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09374_ (.A1(_03993_),
    .A2(_03996_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09375_ (.A1(_04060_),
    .A2(_04053_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09376_ (.A1(_03982_),
    .A2(_03987_),
    .A3(_03988_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09377_ (.A1(_03997_),
    .A2(_03999_),
    .A3(_04062_),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09378_ (.A1(_04051_),
    .A2(_04052_),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09379_ (.A1(_04051_),
    .A2(_04052_),
    .Z(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09380_ (.A1(_04048_),
    .A2(_04064_),
    .B(_04065_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09381_ (.A1(_04061_),
    .A2(_04063_),
    .A3(_04066_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09382_ (.A1(_04067_),
    .A2(_04059_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09383_ (.A1(net354),
    .A2(_04067_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09384_ (.A1(_04057_),
    .A2(_04068_),
    .B(_04069_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09385_ (.A1(_04051_),
    .A2(_04052_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09386_ (.A1(_04048_),
    .A2(_04064_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09387_ (.A1(_04071_),
    .A2(_04072_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09388_ (.A1(_04061_),
    .A2(_04063_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09389_ (.A1(_04061_),
    .A2(_04063_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09390_ (.A1(_04073_),
    .A2(_04074_),
    .B(_04075_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09391_ (.A1(_04002_),
    .A2(_04003_),
    .A3(_03991_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09392_ (.A1(_04076_),
    .A2(_04077_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09393_ (.A1(_04076_),
    .A2(_04077_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09394_ (.A1(_04070_),
    .A2(_04078_),
    .B(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09395_ (.A1(_04006_),
    .A2(_04007_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09396_ (.A1(_03972_),
    .A2(_03980_),
    .B1(_04008_),
    .B2(_04080_),
    .C(_04081_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09397_ (.A1(_03902_),
    .A2(_03906_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09398_ (.A1(_04083_),
    .A2(_03927_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09399_ (.A1(_03977_),
    .A2(_03978_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09400_ (.A1(_03973_),
    .A2(_03979_),
    .B(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09401_ (.A1(_04084_),
    .A2(_04086_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09402_ (.A1(_04084_),
    .A2(_04086_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09403_ (.A1(_03981_),
    .A2(_04082_),
    .A3(_04087_),
    .B(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09404_ (.A1(_03912_),
    .A2(_03925_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09405_ (.A1(_03910_),
    .A2(_03926_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09406_ (.A1(_03919_),
    .A2(_03923_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09407_ (.A1(_03916_),
    .A2(_03924_),
    .B(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09408_ (.A1(_00730_),
    .A2(_01012_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09409_ (.A1(_00758_),
    .A2(_01030_),
    .B1(_00827_),
    .B2(_00720_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09410_ (.A1(_00719_),
    .A2(_00757_),
    .A3(_01030_),
    .A4(_00827_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09411_ (.A1(_03922_),
    .A2(_04095_),
    .B(_04096_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09412_ (.I(_04097_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09413_ (.A1(_00775_),
    .A2(_00793_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09414_ (.A1(_00718_),
    .A2(_03892_),
    .A3(_03888_),
    .A4(_01028_),
    .Z(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09415_ (.A1(_00757_),
    .A2(_03888_),
    .B1(_01029_),
    .B2(_00719_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09416_ (.A1(_04100_),
    .A2(_04101_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09417_ (.A1(_04099_),
    .A2(_04102_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09418_ (.A1(_04098_),
    .A2(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09419_ (.A1(_04094_),
    .A2(_04104_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09420_ (.A1(_04093_),
    .A2(_04105_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09421_ (.A1(_03915_),
    .A2(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09422_ (.A1(_04090_),
    .A2(_04091_),
    .B(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09423_ (.A1(_04099_),
    .A2(_04102_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09424_ (.A1(_00764_),
    .A2(_00774_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09425_ (.A1(_00720_),
    .A2(_01024_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09426_ (.A1(_00730_),
    .A2(_00793_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09427_ (.A1(_04110_),
    .A2(_04111_),
    .A3(_04112_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09428_ (.A1(_04100_),
    .A2(_04109_),
    .B(_04113_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09429_ (.I(_04114_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09430_ (.A1(_04100_),
    .A2(_04109_),
    .A3(_04113_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09431_ (.A1(_04115_),
    .A2(_04116_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09432_ (.A1(net218),
    .A2(net191),
    .A3(_04104_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09433_ (.A1(_04098_),
    .A2(_04103_),
    .B(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09434_ (.A1(_04117_),
    .A2(_04119_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09435_ (.A1(_04093_),
    .A2(_04105_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09436_ (.A1(_03915_),
    .A2(_04106_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09437_ (.A1(_04121_),
    .A2(_04122_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09438_ (.A1(_04120_),
    .A2(_04123_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09439_ (.A1(_04108_),
    .A2(_04124_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09440_ (.A1(_04090_),
    .A2(_04091_),
    .A3(_04107_),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09441_ (.A1(_04108_),
    .A2(_04126_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09442_ (.A1(_03928_),
    .A2(_04089_),
    .B(_04125_),
    .C(_04127_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09443_ (.A1(_04121_),
    .A2(_04122_),
    .B(_04120_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09444_ (.A1(_04108_),
    .A2(_04124_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09445_ (.A1(_04129_),
    .A2(_04130_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09446_ (.I(_04110_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09447_ (.A1(_00721_),
    .A2(_01025_),
    .B(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09448_ (.A1(net194),
    .A2(_01025_),
    .A3(_04132_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09449_ (.A1(_04133_),
    .A2(_04112_),
    .B(_04134_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09450_ (.A1(_00721_),
    .A2(_00767_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09451_ (.A1(net218),
    .A2(net193),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09452_ (.A1(_04136_),
    .A2(_04137_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09453_ (.I(_04138_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09454_ (.A1(_04135_),
    .A2(_04139_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09455_ (.A1(_04117_),
    .A2(_04119_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09456_ (.A1(_04115_),
    .A2(_04141_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09457_ (.A1(_04140_),
    .A2(_04142_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09458_ (.A1(_04128_),
    .A2(_04131_),
    .B(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09459_ (.A1(_04140_),
    .A2(_04141_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09460_ (.I(_04145_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09461_ (.A1(_04135_),
    .A2(_04139_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09462_ (.A1(_04140_),
    .A2(_04115_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09463_ (.A1(_04147_),
    .A2(_04148_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09464_ (.A1(_00727_),
    .A2(_00722_),
    .A3(_04132_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09465_ (.A1(_04149_),
    .A2(_04150_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09466_ (.A1(_04146_),
    .A2(_04151_),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09467_ (.A1(_04146_),
    .A2(_04151_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09468_ (.A1(_04132_),
    .A2(_04149_),
    .B(net218),
    .C(net194),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09469_ (.A1(_04153_),
    .A2(_04154_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09470_ (.A1(_04144_),
    .A2(_04152_),
    .B(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09471_ (.A1(_04144_),
    .A2(_04152_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09472_ (.A1(_04143_),
    .A2(_04128_),
    .A3(_04131_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09473_ (.A1(_04144_),
    .A2(_04158_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09474_ (.A1(_04127_),
    .A2(_03928_),
    .A3(_04089_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09475_ (.A1(_03928_),
    .A2(_04089_),
    .B(_04127_),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09476_ (.A1(_04125_),
    .A2(_04161_),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09477_ (.A1(_03981_),
    .A2(_04082_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09478_ (.A1(_04084_),
    .A2(_04086_),
    .A3(_04163_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09479_ (.A1(_04008_),
    .A2(_04080_),
    .B(_04081_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09480_ (.A1(_03972_),
    .A2(_03980_),
    .A3(_04165_),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09481_ (.A1(_04008_),
    .A2(_04080_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09482_ (.A1(_04070_),
    .A2(_04078_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09483_ (.A1(_04057_),
    .A2(_04068_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(_04025_),
    .A2(_04043_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09485_ (.A1(_04170_),
    .A2(_04056_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09486_ (.A1(_04032_),
    .A2(_04041_),
    .A3(_04042_),
    .Z(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09487_ (.A1(_04043_),
    .A2(_04172_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09488_ (.A1(_04039_),
    .A2(_04040_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09489_ (.A1(_04035_),
    .A2(_04038_),
    .Z(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(_04036_),
    .A2(_04037_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09491_ (.A1(_01491_),
    .A2(_01021_),
    .B(_04175_),
    .C(_04176_),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09492_ (.A1(_04171_),
    .A2(_04173_),
    .A3(_04174_),
    .A4(_04177_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09493_ (.A1(_04168_),
    .A2(_04169_),
    .A3(_04178_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09494_ (.A1(_04164_),
    .A2(_04166_),
    .A3(_04167_),
    .A4(_04179_),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09495_ (.A1(_04160_),
    .A2(_04162_),
    .A3(_04180_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _09496_ (.A1(_04157_),
    .A2(_04159_),
    .A3(_04181_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09497_ (.A1(_01229_),
    .A2(_01285_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09498_ (.A1(_04156_),
    .A2(_04182_),
    .B(_04183_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09499_ (.A1(_01129_),
    .A2(_03587_),
    .A3(_01511_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09500_ (.I(_04185_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09501_ (.A1(_01575_),
    .A2(_01578_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09502_ (.A1(_01510_),
    .A2(_03151_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09503_ (.A1(_04187_),
    .A2(_04188_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09504_ (.A1(_03736_),
    .A2(_03416_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09505_ (.A1(_04189_),
    .A2(_04190_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09506_ (.A1(\as2650.debug_psl[6] ),
    .A2(_02477_),
    .B(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09507_ (.A1(_01856_),
    .A2(_04186_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09508_ (.I(_00833_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09509_ (.A1(net217),
    .A2(net216),
    .A3(net215),
    .A4(_01492_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09510_ (.A1(_04194_),
    .A2(_01768_),
    .A3(_01747_),
    .A4(_04195_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09511_ (.A1(_04184_),
    .A2(_04186_),
    .A3(_04192_),
    .B1(_04193_),
    .B2(_04196_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09512_ (.A1(_03834_),
    .A2(_03835_),
    .B(_03824_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09513_ (.A1(_03607_),
    .A2(_03647_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09514_ (.A1(_04198_),
    .A2(_04199_),
    .B(_03683_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09515_ (.A1(_03686_),
    .A2(_03650_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09516_ (.A1(_03653_),
    .A2(_03688_),
    .B1(_04200_),
    .B2(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09517_ (.A1(_03689_),
    .A2(_03685_),
    .A3(_03687_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09518_ (.A1(_03689_),
    .A2(_03652_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09519_ (.I(_03653_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09520_ (.A1(_01703_),
    .A2(_04205_),
    .B(_03688_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09521_ (.A1(_03689_),
    .A2(_03841_),
    .B1(_04206_),
    .B2(_02920_),
    .C(_03842_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09522_ (.A1(_01168_),
    .A2(_04204_),
    .B(_04207_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09523_ (.A1(_01200_),
    .A2(_04202_),
    .A3(_04203_),
    .B(_04208_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09524_ (.A1(_03594_),
    .A2(_03842_),
    .B(_04209_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09525_ (.A1(_03683_),
    .A2(_03649_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09526_ (.A1(_03684_),
    .A2(_03680_),
    .A3(_03681_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09527_ (.A1(_03823_),
    .A2(_04200_),
    .A3(_04212_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09528_ (.A1(_01283_),
    .A2(_03682_),
    .B(_03603_),
    .C(_02920_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09529_ (.A1(_03684_),
    .A2(_03773_),
    .B1(_03776_),
    .B2(_03600_),
    .C(_04214_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09530_ (.A1(_02469_),
    .A2(_04211_),
    .B(_04213_),
    .C(_04215_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09531_ (.A1(_03622_),
    .A2(_03639_),
    .B(_03644_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09532_ (.A1(_03833_),
    .A2(_04217_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09533_ (.A1(_03833_),
    .A2(_03831_),
    .A3(_03832_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09534_ (.A1(_03613_),
    .A2(_03615_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09535_ (.A1(_02467_),
    .A2(_04220_),
    .B(_03675_),
    .C(_02564_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09536_ (.A1(_03676_),
    .A2(_03772_),
    .B1(_03775_),
    .B2(_03613_),
    .C(_04221_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09537_ (.A1(_01200_),
    .A2(_03677_),
    .A3(_04219_),
    .B(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09538_ (.A1(_01168_),
    .A2(_04218_),
    .B(_04223_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09539_ (.A1(_03672_),
    .A2(_03668_),
    .A3(_03669_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09540_ (.A1(_01199_),
    .A2(_03831_),
    .A3(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09541_ (.A1(_03672_),
    .A2(_03639_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09542_ (.A1(_03619_),
    .A2(_03671_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09543_ (.A1(_02565_),
    .A2(_04228_),
    .B1(_03726_),
    .B2(_03644_),
    .C(_03774_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09544_ (.A1(_03672_),
    .A2(_03841_),
    .B1(_04227_),
    .B2(_02468_),
    .C(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _09545_ (.A1(_03670_),
    .A2(_03842_),
    .B1(_04226_),
    .B2(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09546_ (.A1(_03635_),
    .A2(_03662_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09547_ (.A1(_04232_),
    .A2(_03634_),
    .B(_02468_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09548_ (.A1(_04232_),
    .A2(_03634_),
    .B(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09549_ (.A1(_04232_),
    .A2(_03826_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09550_ (.A1(_03823_),
    .A2(_03664_),
    .A3(_04235_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09551_ (.A1(_01703_),
    .A2(_03635_),
    .B(_03632_),
    .C(_01231_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09552_ (.A1(_04232_),
    .A2(_03773_),
    .B1(_03775_),
    .B2(_03661_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09553_ (.A1(_04234_),
    .A2(_04236_),
    .A3(_04237_),
    .A4(_04238_),
    .Z(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09554_ (.A1(_03627_),
    .A2(_03636_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09555_ (.A1(_03667_),
    .A2(_03664_),
    .A3(_03665_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09556_ (.A1(_03822_),
    .A2(_03829_),
    .A3(_04241_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09557_ (.A1(_01282_),
    .A2(_03638_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09558_ (.A1(_03637_),
    .A2(_03666_),
    .B(_04243_),
    .C(_01231_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09559_ (.A1(_03667_),
    .A2(_03773_),
    .B1(_03775_),
    .B2(_03637_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09560_ (.A1(_04242_),
    .A2(_04244_),
    .A3(_04245_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09561_ (.A1(_01168_),
    .A2(_04240_),
    .B(_04246_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09562_ (.A1(_04224_),
    .A2(_04231_),
    .A3(_04239_),
    .A4(_04247_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09563_ (.A1(_03847_),
    .A2(_04248_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09564_ (.A1(_04216_),
    .A2(_04249_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09565_ (.A1(_03780_),
    .A2(_03781_),
    .B1(_04210_),
    .B2(_04250_),
    .C(_03724_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09566_ (.A1(_03160_),
    .A2(_03768_),
    .B1(_03725_),
    .B2(_04197_),
    .C(_04251_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09567_ (.A1(_01855_),
    .A2(_03744_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09568_ (.A1(_01026_),
    .A2(_01656_),
    .B1(net215),
    .B2(_01388_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09569_ (.A1(_01031_),
    .A2(_01388_),
    .B1(_01501_),
    .B2(_01390_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09570_ (.A1(_04194_),
    .A2(_01401_),
    .B1(_01768_),
    .B2(_01349_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09571_ (.A1(_01497_),
    .A2(_01614_),
    .B1(_01491_),
    .B2(_01598_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(_01497_),
    .A2(_01353_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09573_ (.A1(net210),
    .A2(_01625_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09574_ (.A1(_04257_),
    .A2(_04258_),
    .B(_04259_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09575_ (.A1(_04256_),
    .A2(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09576_ (.A1(_04255_),
    .A2(_04261_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09577_ (.A1(_01026_),
    .A2(_01656_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09578_ (.A1(_04254_),
    .A2(_04262_),
    .B(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09579_ (.A1(net217),
    .A2(_01418_),
    .B(_04264_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09580_ (.A1(_01855_),
    .A2(_03744_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09581_ (.A1(_01667_),
    .A2(_03855_),
    .B(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09582_ (.A1(_04253_),
    .A2(_04267_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09583_ (.A1(\as2650.debug_psl[1] ),
    .A2(_04266_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09584_ (.A1(\as2650.debug_psl[1] ),
    .A2(_04253_),
    .B1(_04265_),
    .B2(_04268_),
    .C(_04269_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09585_ (.A1(net199),
    .A2(_01615_),
    .B1(_01492_),
    .B2(_01598_),
    .C(_04267_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09586_ (.A1(_04255_),
    .A2(_04256_),
    .A3(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09587_ (.A1(_03658_),
    .A2(_03741_),
    .B(_04258_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09588_ (.A1(_01837_),
    .A2(_03856_),
    .B(_04253_),
    .C(_04254_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09589_ (.A1(_04263_),
    .A2(_04259_),
    .A3(_04273_),
    .A4(_04274_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09590_ (.A1(_04272_),
    .A2(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09591_ (.A1(_03160_),
    .A2(_03768_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09592_ (.A1(_04270_),
    .A2(_04276_),
    .B(_04277_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09593_ (.A1(_01779_),
    .A2(_01599_),
    .B(_03633_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09594_ (.I(_04279_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09595_ (.A1(_03728_),
    .A2(_04280_),
    .B(_03730_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09596_ (.I(_01383_),
    .Z(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09597_ (.A1(_01637_),
    .A2(_01625_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09598_ (.A1(_01674_),
    .A2(_01418_),
    .A3(_01648_),
    .A4(_01615_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09599_ (.A1(_04282_),
    .A2(_03731_),
    .A3(_04283_),
    .A4(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09600_ (.A1(_03728_),
    .A2(_04252_),
    .A3(_04278_),
    .B1(_04281_),
    .B2(_04285_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09601_ (.A1(_03732_),
    .A2(_03745_),
    .B(_03663_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09602_ (.A1(_01361_),
    .A2(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09603_ (.A1(_01664_),
    .A2(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09604_ (.A1(_03731_),
    .A2(_04289_),
    .B(_03721_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09605_ (.A1(_02665_),
    .A2(_02470_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09606_ (.A1(_02579_),
    .A2(_01837_),
    .A3(_02471_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09607_ (.A1(_04286_),
    .A2(_04290_),
    .B(_04291_),
    .C(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _09608_ (.A1(\as2650.debug_psu[5] ),
    .A2(\as2650.debug_psu[4] ),
    .A3(net306),
    .A4(_02546_),
    .Z(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09609_ (.A1(\as2650.debug_psu[7] ),
    .A2(_02465_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09610_ (.A1(_01754_),
    .A2(\as2650.debug_psl[2] ),
    .A3(_03732_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09611_ (.A1(_01806_),
    .A2(_01559_),
    .A3(_03580_),
    .A4(_01568_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09612_ (.A1(_04296_),
    .A2(_04297_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09613_ (.A1(_01564_),
    .A2(_03720_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09614_ (.A1(_01576_),
    .A2(_02470_),
    .Z(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09615_ (.A1(_04294_),
    .A2(_04295_),
    .B1(_04298_),
    .B2(_04299_),
    .C(_04300_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09616_ (.A1(_02943_),
    .A2(_04301_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09617_ (.A1(_01429_),
    .A2(_01201_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09618_ (.A1(_01559_),
    .A2(_02943_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09619_ (.A1(_04293_),
    .A2(_04302_),
    .B(_04303_),
    .C(_04304_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09620_ (.A1(_01092_),
    .A2(_03720_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09621_ (.I(_01577_),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09622_ (.A1(_01568_),
    .A2(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09623_ (.A1(_02576_),
    .A2(_04306_),
    .A3(_04308_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09624_ (.A1(_03732_),
    .A2(_04307_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09625_ (.A1(_01923_),
    .A2(_02466_),
    .B(_02619_),
    .C(_04310_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09626_ (.A1(_04309_),
    .A2(_04311_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09627_ (.A1(_04295_),
    .A2(_04299_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09628_ (.A1(_01682_),
    .A2(_03720_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09629_ (.A1(_01771_),
    .A2(_04307_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09630_ (.A1(_02615_),
    .A2(_04314_),
    .A3(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09631_ (.A1(_02813_),
    .A2(_04313_),
    .B(_04316_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09632_ (.I0(_01754_),
    .I1(_01886_),
    .S(_02578_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09633_ (.A1(_01872_),
    .A2(_00687_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09634_ (.A1(_01558_),
    .A2(_00687_),
    .B(_04319_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09635_ (.A1(_01950_),
    .A2(_01577_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09636_ (.A1(_01559_),
    .A2(_02465_),
    .B(_04321_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09637_ (.A1(\as2650.debug_psu[4] ),
    .A2(_02578_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09638_ (.A1(_01806_),
    .A2(_02465_),
    .B(_04323_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09639_ (.A1(_02801_),
    .A2(_04322_),
    .B1(_04324_),
    .B2(_02626_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09640_ (.A1(_02676_),
    .A2(_04318_),
    .B1(_04320_),
    .B2(_02658_),
    .C(_04325_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09641_ (.A1(_04303_),
    .A2(_04312_),
    .A3(_04317_),
    .A4(_04326_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09642_ (.A1(_03717_),
    .A2(_04327_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09643_ (.A1(_03159_),
    .A2(_02802_),
    .A3(_03707_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09644_ (.A1(_01560_),
    .A2(_02790_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09645_ (.A1(_04329_),
    .A2(_04330_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09646_ (.A1(_04305_),
    .A2(_04328_),
    .B1(_04331_),
    .B2(_03717_),
    .C(_03769_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09647_ (.A1(_02812_),
    .A2(_01677_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09648_ (.A1(_02813_),
    .A2(_01677_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09649_ (.A1(_02827_),
    .A2(_01669_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09650_ (.A1(_02827_),
    .A2(_01669_),
    .B(_04333_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09651_ (.A1(_04334_),
    .A2(_04336_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09652_ (.A1(_02769_),
    .A2(_01660_),
    .B(_04335_),
    .C(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09653_ (.A1(_02765_),
    .A2(_01651_),
    .B1(_01660_),
    .B2(_02769_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09654_ (.A1(_02765_),
    .A2(_01651_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09655_ (.A1(_02726_),
    .A2(_01643_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09656_ (.A1(_04340_),
    .A2(_04341_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09657_ (.A1(_02645_),
    .A2(_01608_),
    .B1(_01632_),
    .B2(_02715_),
    .C1(_01621_),
    .C2(_02675_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09658_ (.A1(_02715_),
    .A2(_01632_),
    .B(_01621_),
    .C(_02675_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09659_ (.A1(_02715_),
    .A2(_01632_),
    .B1(_01643_),
    .B2(_02726_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09660_ (.A1(_04343_),
    .A2(_04344_),
    .A3(_04345_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09661_ (.A1(_04342_),
    .A2(_04346_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09662_ (.A1(_04339_),
    .A2(_04347_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09663_ (.A1(_04334_),
    .A2(_04335_),
    .B1(_04338_),
    .B2(_04348_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09664_ (.A1(\as2650.debug_psl[1] ),
    .A2(_04334_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09665_ (.A1(_01754_),
    .A2(_04333_),
    .B(_04350_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09666_ (.A1(_04333_),
    .A2(_04349_),
    .B(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09667_ (.A1(_03768_),
    .A2(_04352_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09668_ (.A1(_01749_),
    .A2(_01191_),
    .A3(_01342_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09669_ (.A1(_04353_),
    .A2(_04354_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09670_ (.A1(_02676_),
    .A2(_01372_),
    .B1(_03741_),
    .B2(_02658_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09671_ (.A1(_03745_),
    .A2(_02814_),
    .B1(_02790_),
    .B2(_03857_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09672_ (.I(_01349_),
    .Z(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09673_ (.A1(_04358_),
    .A2(_02716_),
    .B1(_02766_),
    .B2(_03858_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09674_ (.I(_01401_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09675_ (.A1(_04360_),
    .A2(_02731_),
    .B1(_02770_),
    .B2(_04282_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09676_ (.A1(_04356_),
    .A2(_04357_),
    .A3(_04359_),
    .A4(_04361_),
    .Z(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09677_ (.A1(_04332_),
    .A2(_04355_),
    .B1(_04362_),
    .B2(_04354_),
    .C(_03699_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _09678_ (.I(_04210_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09679_ (.I(_03783_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09680_ (.A1(_04364_),
    .A2(_04216_),
    .A3(_04249_),
    .B(_04365_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09681_ (.A1(_03716_),
    .A2(_04366_),
    .B(_02562_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09682_ (.A1(_02583_),
    .A2(_03699_),
    .B(_03799_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09683_ (.A1(_04293_),
    .A2(_04302_),
    .B(_04304_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09684_ (.A1(_02562_),
    .A2(_04369_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09685_ (.A1(_04363_),
    .A2(_04367_),
    .B(_04368_),
    .C(_04370_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09686_ (.A1(\as2650.cycle[8] ),
    .A2(_01539_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09687_ (.I(_04372_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09688_ (.A1(_03716_),
    .A2(_04366_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09689_ (.A1(_04353_),
    .A2(_04374_),
    .B(_03799_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09690_ (.A1(_04373_),
    .A2(_04375_),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09691_ (.A1(_02607_),
    .A2(_02640_),
    .A3(_02616_),
    .A4(_02619_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09692_ (.A1(_02766_),
    .A2(_02791_),
    .A3(_02781_),
    .A4(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09693_ (.A1(_02814_),
    .A2(_04373_),
    .A3(_04378_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09694_ (.A1(\as2650.cycle[10] ),
    .A2(_01528_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09695_ (.A1(_04371_),
    .A2(_04376_),
    .B(_04379_),
    .C(_04380_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09696_ (.I0(net2),
    .I1(net26),
    .I2(net10),
    .I3(net18),
    .S0(\as2650.ext_io_addr[6] ),
    .S1(_01518_),
    .Z(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09697_ (.I(\as2650.ext_io_addr[7] ),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09698_ (.I(\as2650.ext_io_addr[6] ),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09699_ (.I0(net3),
    .I1(net11),
    .I2(net27),
    .I3(net19),
    .S0(_04383_),
    .S1(_04384_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09700_ (.I0(net5),
    .I1(net13),
    .I2(net29),
    .I3(net21),
    .S0(_01518_),
    .S1(_01520_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _09701_ (.I0(net1),
    .I1(net9),
    .I2(net25),
    .I3(net17),
    .S0(_04383_),
    .S1(_04384_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _09702_ (.I0(net6),
    .I1(net30),
    .I2(net14),
    .I3(net22),
    .S0(\as2650.ext_io_addr[6] ),
    .S1(_01518_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09703_ (.I0(net7),
    .I1(net15),
    .I2(net31),
    .I3(net23),
    .S0(_04383_),
    .S1(_04384_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09704_ (.I0(net4),
    .I1(net12),
    .I2(net28),
    .I3(net20),
    .S0(_04383_),
    .S1(_01520_),
    .Z(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09705_ (.A1(_04387_),
    .A2(_04388_),
    .A3(_04389_),
    .A4(_04390_),
    .Z(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09706_ (.A1(_04382_),
    .A2(_04385_),
    .A3(_04386_),
    .A4(_04391_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09707_ (.I0(net8),
    .I1(net16),
    .I2(net32),
    .I3(net24),
    .S0(\as2650.ext_io_addr[7] ),
    .S1(_04384_),
    .Z(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09708_ (.A1(_04392_),
    .A2(_04393_),
    .B(_01477_),
    .C(_01529_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09709_ (.A1(_02670_),
    .A2(_04381_),
    .A3(_04394_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09710_ (.I(_04395_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09711_ (.A1(_02658_),
    .A2(_01608_),
    .B1(_01621_),
    .B2(_02676_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09712_ (.A1(_04339_),
    .A2(_04342_),
    .A3(_04345_),
    .A4(_04396_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09713_ (.A1(_04338_),
    .A2(_04343_),
    .A3(_04397_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09714_ (.A1(_04352_),
    .A2(_04398_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09715_ (.I(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09716_ (.A1(_02587_),
    .A2(_04365_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09717_ (.A1(_03769_),
    .A2(_04400_),
    .B(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09718_ (.A1(_03799_),
    .A2(_04402_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09719_ (.A1(_02590_),
    .A2(_02567_),
    .B(_02991_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09720_ (.A1(_01564_),
    .A2(_02991_),
    .B(_03718_),
    .C(_04404_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09721_ (.A1(_02583_),
    .A2(_04400_),
    .B(_04354_),
    .C(_02586_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09722_ (.A1(_02583_),
    .A2(_04405_),
    .B(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09723_ (.A1(_04401_),
    .A2(_04407_),
    .B(_03703_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09724_ (.I(_04270_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09725_ (.A1(_01564_),
    .A2(_03736_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09726_ (.A1(_02477_),
    .A2(_03440_),
    .B(_04189_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09727_ (.A1(_04183_),
    .A2(_04156_),
    .B1(_04410_),
    .B2(_04411_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09728_ (.A1(_04186_),
    .A2(_04412_),
    .B(_04193_),
    .C(_03724_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09729_ (.A1(_03729_),
    .A2(_02585_),
    .A3(_03782_),
    .B(_04413_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09730_ (.I0(_04409_),
    .I1(_04414_),
    .S(_04277_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09731_ (.A1(_03728_),
    .A2(_04415_),
    .B(_04281_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09732_ (.A1(_03857_),
    .A2(_03731_),
    .B(_03721_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09733_ (.A1(_01856_),
    .A2(_03722_),
    .B1(_04416_),
    .B2(_04417_),
    .C(_04291_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09734_ (.A1(_04291_),
    .A2(_04313_),
    .B(_04418_),
    .C(_02944_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09735_ (.A1(_03709_),
    .A2(_01201_),
    .B(_03717_),
    .C(_04406_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09736_ (.A1(_01565_),
    .A2(_03714_),
    .B1(_04420_),
    .B2(_02562_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09737_ (.A1(_04419_),
    .A2(_04421_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09738_ (.A1(_04408_),
    .A2(_04422_),
    .B(_04368_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09739_ (.A1(_04403_),
    .A2(_04423_),
    .B(_04372_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09740_ (.A1(_02813_),
    .A2(_04372_),
    .B(_04380_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09741_ (.I(_04425_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09742_ (.A1(_04380_),
    .A2(_04393_),
    .B(_03182_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09743_ (.A1(_04424_),
    .A2(_04426_),
    .B(_04427_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09744_ (.I(_01087_),
    .Z(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09745_ (.A1(_01261_),
    .A2(_01324_),
    .A3(_01705_),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09746_ (.A1(_02559_),
    .A2(_02568_),
    .B(_02560_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09747_ (.A1(_02560_),
    .A2(_04429_),
    .B(_04430_),
    .C(_01453_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09748_ (.I(_03735_),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09749_ (.A1(_01700_),
    .A2(_04432_),
    .A3(_02557_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09750_ (.A1(_01874_),
    .A2(_04433_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09751_ (.A1(_02484_),
    .A2(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09752_ (.A1(net188),
    .A2(_02473_),
    .B(_04435_),
    .C(_01275_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09753_ (.A1(_01874_),
    .A2(_01102_),
    .B(_04436_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09754_ (.A1(_04431_),
    .A2(_04437_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09755_ (.I(_02588_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09756_ (.I(_01872_),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09757_ (.A1(_04440_),
    .A2(_02640_),
    .B(_03708_),
    .C(_03710_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09758_ (.A1(_02708_),
    .A2(_04439_),
    .A3(_04441_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09759_ (.I(_01704_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09760_ (.A1(_04443_),
    .A2(_02666_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09761_ (.I(_04444_),
    .Z(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09762_ (.A1(_04438_),
    .A2(_04442_),
    .B(_04445_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09763_ (.A1(_02666_),
    .A2(_03065_),
    .B(_04440_),
    .C(_04443_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09764_ (.A1(_04446_),
    .A2(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09765_ (.A1(_04428_),
    .A2(_04448_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09766_ (.I(_02472_),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09767_ (.A1(_03141_),
    .A2(_03143_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09768_ (.A1(_04432_),
    .A2(_02556_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09769_ (.A1(_04440_),
    .A2(_01701_),
    .B(_04451_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09770_ (.A1(_04450_),
    .A2(_04452_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09771_ (.A1(_02473_),
    .A2(_04453_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09772_ (.A1(net199),
    .A2(_04449_),
    .B(_04454_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09773_ (.A1(_01887_),
    .A2(_02599_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09774_ (.A1(_02599_),
    .A2(_04455_),
    .B(_04456_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09775_ (.A1(_01887_),
    .A2(_02607_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09776_ (.A1(_01268_),
    .A2(_04450_),
    .A3(_04429_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09777_ (.A1(_04439_),
    .A2(_03761_),
    .A3(_04458_),
    .B(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09778_ (.A1(_04431_),
    .A2(_04457_),
    .B1(_04460_),
    .B2(_01454_),
    .C(_04445_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09779_ (.A1(_04443_),
    .A2(_04450_),
    .A3(_03128_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09780_ (.A1(_01526_),
    .A2(_04461_),
    .A3(_04462_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09781_ (.A1(_01902_),
    .A2(_01288_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09782_ (.I(_04451_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09783_ (.A1(_01682_),
    .A2(_03514_),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09784_ (.I0(_04465_),
    .I1(_01901_),
    .S(_01701_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09785_ (.A1(_04464_),
    .A2(_04466_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09786_ (.A1(_02521_),
    .A2(_04464_),
    .B(_04467_),
    .C(_02484_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09787_ (.A1(net210),
    .A2(_04449_),
    .B(_04468_),
    .C(_02598_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09788_ (.A1(_04463_),
    .A2(_04469_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09789_ (.A1(_01902_),
    .A2(_02617_),
    .B(_03794_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09790_ (.A1(_01316_),
    .A2(_04429_),
    .A3(_04465_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09791_ (.A1(_04439_),
    .A2(_04471_),
    .B(_04472_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09792_ (.A1(_04431_),
    .A2(_04470_),
    .B1(_04473_),
    .B2(_01454_),
    .C(_04445_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09793_ (.A1(_02573_),
    .A2(_01706_),
    .A3(_04465_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09794_ (.A1(_01526_),
    .A2(_04474_),
    .A3(_04475_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09795_ (.A1(_01681_),
    .A2(_03142_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09796_ (.A1(_01684_),
    .A2(_03143_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09797_ (.A1(_01683_),
    .A2(_04476_),
    .B(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09798_ (.A1(_04429_),
    .A2(_04478_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09799_ (.I(_01683_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09800_ (.A1(_04480_),
    .A2(_02620_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _09801_ (.A1(_03502_),
    .A2(_04443_),
    .A3(_04479_),
    .B1(_04481_),
    .B2(_04439_),
    .B3(_03808_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09802_ (.A1(_01509_),
    .A2(_04476_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09803_ (.A1(_02475_),
    .A2(_04483_),
    .B(_02665_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09804_ (.A1(_01701_),
    .A2(_04477_),
    .B1(_04484_),
    .B2(_04480_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09805_ (.A1(_02557_),
    .A2(_04485_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09806_ (.A1(_02552_),
    .A2(_04464_),
    .B(_04486_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09807_ (.A1(_02484_),
    .A2(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09808_ (.A1(net214),
    .A2(_04449_),
    .B(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09809_ (.I(_04430_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09810_ (.A1(_02560_),
    .A2(_04479_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09811_ (.A1(_01468_),
    .A2(_04490_),
    .A3(_04491_),
    .B1(_02598_),
    .B2(_04480_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09812_ (.A1(_02599_),
    .A2(_04489_),
    .B(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09813_ (.A1(_02748_),
    .A2(_04482_),
    .B(_04493_),
    .C(_04444_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09814_ (.A1(_04445_),
    .A2(_04478_),
    .B(_04494_),
    .C(_03534_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09815_ (.A1(_02473_),
    .A2(_03754_),
    .A3(_03573_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09816_ (.A1(_01804_),
    .A2(_02485_),
    .B(_04495_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09817_ (.A1(_01931_),
    .A2(_02480_),
    .B1(_04496_),
    .B2(_02483_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09818_ (.A1(_01931_),
    .A2(_02628_),
    .B(_02589_),
    .C(_03818_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09819_ (.A1(_02570_),
    .A2(_04497_),
    .B1(_04498_),
    .B2(_03049_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09820_ (.A1(_03105_),
    .A2(_04499_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09821_ (.I(_04500_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09822_ (.I(_04329_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09823_ (.A1(net306),
    .A2(_02791_),
    .B(_04501_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09824_ (.A1(_03755_),
    .A2(_03120_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09825_ (.A1(_01838_),
    .A2(_02485_),
    .B(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09826_ (.A1(net181),
    .A2(_02480_),
    .B1(_04504_),
    .B2(_02483_),
    .C(_02569_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09827_ (.A1(_02570_),
    .A2(_04502_),
    .B(_04505_),
    .C(_03534_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09828_ (.A1(_04449_),
    .A2(_03754_),
    .A3(_03146_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09829_ (.A1(_01857_),
    .A2(_02485_),
    .B(_04506_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09830_ (.A1(net37),
    .A2(_02480_),
    .B1(_04507_),
    .B2(_02483_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09831_ (.A1(\as2650.debug_psu[7] ),
    .A2(_02992_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09832_ (.A1(_02568_),
    .A2(_04509_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09833_ (.A1(_01306_),
    .A2(_02589_),
    .A3(_04404_),
    .A4(_04510_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09834_ (.A1(_02570_),
    .A2(_04508_),
    .B(_04511_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09835_ (.A1(_03105_),
    .A2(_04512_),
    .Z(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09836_ (.I(_04513_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09837_ (.I(_01516_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09838_ (.I0(net44),
    .I1(\as2650.irqs_latch[1] ),
    .S(_04514_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09839_ (.I(_04515_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09840_ (.A1(net45),
    .A2(_00010_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09841_ (.A1(_02693_),
    .A2(_00010_),
    .B(_04516_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09842_ (.I0(net46),
    .I1(\as2650.irqs_latch[3] ),
    .S(_04514_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09843_ (.I(_04517_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09844_ (.I0(\as2650.trap ),
    .I1(\as2650.irqs_latch[4] ),
    .S(_04514_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09845_ (.I(_04518_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09846_ (.I0(net47),
    .I1(\as2650.irqs_latch[5] ),
    .S(_04514_),
    .Z(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09847_ (.I(_04519_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09848_ (.I0(net48),
    .I1(\as2650.irqs_latch[6] ),
    .S(_01516_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09849_ (.I(_04520_),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09850_ (.I0(net49),
    .I1(\as2650.irqs_latch[7] ),
    .S(_01516_),
    .Z(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09851_ (.I(_04521_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09852_ (.I(_02534_),
    .Z(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09853_ (.A1(_01901_),
    .A2(_01924_),
    .Z(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09854_ (.A1(_01961_),
    .A2(_04522_),
    .A3(_04523_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09855_ (.I(_04524_),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09856_ (.I(_04525_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09857_ (.I(_04524_),
    .Z(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09858_ (.I(_04527_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09859_ (.A1(\as2650.stack[5][0] ),
    .A2(_04528_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09860_ (.A1(_01737_),
    .A2(_04526_),
    .B(_04529_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09861_ (.A1(\as2650.stack[5][1] ),
    .A2(_04528_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09862_ (.A1(_01760_),
    .A2(_04526_),
    .B(_04530_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09863_ (.A1(\as2650.stack[5][2] ),
    .A2(_04528_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09864_ (.A1(_01777_),
    .A2(_04526_),
    .B(_04531_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09865_ (.A1(\as2650.stack[5][3] ),
    .A2(_04528_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09866_ (.A1(_01801_),
    .A2(_04526_),
    .B(_04532_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09867_ (.I(_04525_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09868_ (.I(_04527_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09869_ (.A1(\as2650.stack[5][4] ),
    .A2(_04534_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09870_ (.A1(_01820_),
    .A2(_04533_),
    .B(_04535_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09871_ (.A1(\as2650.stack[5][5] ),
    .A2(_04534_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09872_ (.A1(_01835_),
    .A2(_04533_),
    .B(_04536_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09873_ (.A1(\as2650.stack[5][6] ),
    .A2(_04534_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09874_ (.A1(_01853_),
    .A2(_04533_),
    .B(_04537_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09875_ (.A1(\as2650.stack[5][7] ),
    .A2(_04534_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09876_ (.A1(_01869_),
    .A2(_04533_),
    .B(_04538_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09877_ (.I(_04525_),
    .Z(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09878_ (.I(_04527_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09879_ (.A1(\as2650.stack[5][8] ),
    .A2(_04540_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09880_ (.A1(_01883_),
    .A2(_04539_),
    .B(_04541_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09881_ (.A1(\as2650.stack[5][9] ),
    .A2(_04540_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09882_ (.A1(_01899_),
    .A2(_04539_),
    .B(_04542_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09883_ (.A1(\as2650.stack[5][10] ),
    .A2(_04540_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09884_ (.A1(_01913_),
    .A2(_04539_),
    .B(_04543_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09885_ (.A1(\as2650.stack[5][11] ),
    .A2(_04540_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09886_ (.A1(_01928_),
    .A2(_04539_),
    .B(_04544_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09887_ (.I(_04525_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09888_ (.I(_04527_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09889_ (.A1(\as2650.stack[5][12] ),
    .A2(_04546_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09890_ (.A1(_01940_),
    .A2(_04545_),
    .B(_04547_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09891_ (.A1(\as2650.stack[5][13] ),
    .A2(_04546_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09892_ (.A1(_01947_),
    .A2(_04545_),
    .B(_04548_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09893_ (.A1(\as2650.stack[5][14] ),
    .A2(_04546_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09894_ (.A1(_01954_),
    .A2(_04545_),
    .B(_04549_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09895_ (.A1(\as2650.stack[5][15] ),
    .A2(_04546_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09896_ (.A1(_01959_),
    .A2(_04545_),
    .B(_04550_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09897_ (.A1(_03158_),
    .A2(_01285_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09898_ (.A1(_02559_),
    .A2(_03403_),
    .A3(_01228_),
    .A4(_04551_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09899_ (.A1(_03153_),
    .A2(_02475_),
    .A3(_04551_),
    .B1(_04552_),
    .B2(\as2650.trap ),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09900_ (.A1(_04428_),
    .A2(_04553_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09901_ (.I(\as2650.cycle[1] ),
    .Z(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09902_ (.I(_04554_),
    .Z(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09903_ (.I(\as2650.cycle[1] ),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09904_ (.I(_03174_),
    .Z(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09905_ (.A1(_04556_),
    .A2(net147),
    .B(_04557_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09906_ (.A1(_04555_),
    .A2(_01599_),
    .B(_04558_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09907_ (.A1(_04556_),
    .A2(net148),
    .B(_04557_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09908_ (.A1(_04555_),
    .A2(_01616_),
    .B(_04559_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09909_ (.A1(_04556_),
    .A2(net149),
    .B(_04557_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09910_ (.A1(_04555_),
    .A2(_01626_),
    .B(_04560_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09911_ (.A1(_04556_),
    .A2(net150),
    .B(_04557_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09912_ (.A1(_04555_),
    .A2(_01637_),
    .B(_04561_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09913_ (.I(_04554_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09914_ (.I(\as2650.cycle[1] ),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09915_ (.I(_03174_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09916_ (.A1(_04563_),
    .A2(net151),
    .B(_04564_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09917_ (.A1(_04562_),
    .A2(_01648_),
    .B(_04565_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09918_ (.A1(_04563_),
    .A2(net152),
    .B(_04564_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09919_ (.A1(_04562_),
    .A2(_01657_),
    .B(_04566_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09920_ (.A1(_04563_),
    .A2(net153),
    .B(_04564_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09921_ (.A1(_04562_),
    .A2(_01664_),
    .B(_04567_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09922_ (.A1(_04563_),
    .A2(net154),
    .B(_04564_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09923_ (.A1(_04562_),
    .A2(_01674_),
    .B(_04568_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09924_ (.A1(_01313_),
    .A2(net146),
    .B(\as2650.cycle[7] ),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09925_ (.A1(_01477_),
    .A2(_04428_),
    .A3(_04569_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09926_ (.I(_01465_),
    .Z(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09927_ (.I(_01546_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09928_ (.I(_04571_),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09929_ (.A1(net140),
    .A2(_01466_),
    .B(_04572_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09930_ (.A1(_02659_),
    .A2(_04570_),
    .B(_04573_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09931_ (.A1(net141),
    .A2(_01466_),
    .B(_04572_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09932_ (.A1(_02677_),
    .A2(_04570_),
    .B(_04574_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09933_ (.A1(net142),
    .A2(_01466_),
    .B(_04572_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09934_ (.A1(_02716_),
    .A2(_04570_),
    .B(_04575_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09935_ (.I(_01464_),
    .Z(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09936_ (.A1(net143),
    .A2(_04576_),
    .B(_04572_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09937_ (.A1(_02739_),
    .A2(_04570_),
    .B(_04577_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09938_ (.I(_01465_),
    .Z(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09939_ (.I(_04571_),
    .Z(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09940_ (.A1(net144),
    .A2(_04576_),
    .B(_04579_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09941_ (.A1(_02766_),
    .A2(_04578_),
    .B(_04580_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09942_ (.A1(net145),
    .A2(_04576_),
    .B(_04579_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09943_ (.A1(_02781_),
    .A2(_04578_),
    .B(_04581_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09944_ (.A1(_01520_),
    .A2(_04576_),
    .B(_04579_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09945_ (.A1(_02791_),
    .A2(_04578_),
    .B(_04582_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09946_ (.A1(_01519_),
    .A2(_01465_),
    .B(_04579_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09947_ (.A1(_02814_),
    .A2(_04578_),
    .B(_04583_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09948_ (.A1(_04554_),
    .A2(_01529_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09949_ (.A1(\as2650.io_bus_we ),
    .A2(_04554_),
    .B(_04584_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09950_ (.A1(_01477_),
    .A2(_04428_),
    .A3(_04585_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09951_ (.I(_01544_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09952_ (.A1(net235),
    .A2(_04586_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09953_ (.A1(_01603_),
    .A2(_04587_),
    .B(_03051_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09954_ (.A1(_00980_),
    .A2(net237),
    .B(_03105_),
    .C(_01618_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09955_ (.A1(net222),
    .A2(_04586_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09956_ (.A1(_01629_),
    .A2(_04588_),
    .B(_03051_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09957_ (.A1(net223),
    .A2(_01545_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09958_ (.A1(_01488_),
    .A2(_01639_),
    .A3(_04589_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09959_ (.A1(net224),
    .A2(_04586_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09960_ (.A1(_01649_),
    .A2(_04590_),
    .B(_01088_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09961_ (.A1(net225),
    .A2(_01545_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09962_ (.A1(_01488_),
    .A2(_01658_),
    .A3(_04591_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09963_ (.A1(net226),
    .A2(_04586_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09964_ (.A1(_01665_),
    .A2(_04592_),
    .B(_01088_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09965_ (.A1(net227),
    .A2(_01545_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09966_ (.A1(_01488_),
    .A2(_01675_),
    .A3(_04593_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09967_ (.A1(_01694_),
    .A2(_01713_),
    .A3(_04523_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09968_ (.I(_04594_),
    .Z(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09969_ (.I(_04595_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09970_ (.I(_04594_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09971_ (.I(_04597_),
    .Z(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09972_ (.A1(\as2650.stack[4][0] ),
    .A2(_04598_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09973_ (.A1(_01737_),
    .A2(_04596_),
    .B(_04599_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09974_ (.A1(\as2650.stack[4][1] ),
    .A2(_04598_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09975_ (.A1(_01760_),
    .A2(_04596_),
    .B(_04600_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09976_ (.A1(\as2650.stack[4][2] ),
    .A2(_04598_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09977_ (.A1(_01777_),
    .A2(_04596_),
    .B(_04601_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09978_ (.A1(\as2650.stack[4][3] ),
    .A2(_04598_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09979_ (.A1(_01801_),
    .A2(_04596_),
    .B(_04602_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09980_ (.I(_04595_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09981_ (.I(_04597_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09982_ (.A1(\as2650.stack[4][4] ),
    .A2(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09983_ (.A1(_01820_),
    .A2(_04603_),
    .B(_04605_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09984_ (.A1(\as2650.stack[4][5] ),
    .A2(_04604_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09985_ (.A1(_01835_),
    .A2(_04603_),
    .B(_04606_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09986_ (.A1(\as2650.stack[4][6] ),
    .A2(_04604_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09987_ (.A1(_01853_),
    .A2(_04603_),
    .B(_04607_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09988_ (.A1(\as2650.stack[4][7] ),
    .A2(_04604_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09989_ (.A1(_01869_),
    .A2(_04603_),
    .B(_04608_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09990_ (.I(_04595_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09991_ (.I(_04597_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09992_ (.A1(\as2650.stack[4][8] ),
    .A2(_04610_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09993_ (.A1(_01883_),
    .A2(_04609_),
    .B(_04611_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09994_ (.A1(\as2650.stack[4][9] ),
    .A2(_04610_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09995_ (.A1(_01899_),
    .A2(_04609_),
    .B(_04612_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09996_ (.A1(\as2650.stack[4][10] ),
    .A2(_04610_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09997_ (.A1(_01913_),
    .A2(_04609_),
    .B(_04613_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09998_ (.A1(\as2650.stack[4][11] ),
    .A2(_04610_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09999_ (.A1(_01928_),
    .A2(_04609_),
    .B(_04614_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10000_ (.I(_04595_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10001_ (.I(_04597_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10002_ (.A1(\as2650.stack[4][12] ),
    .A2(_04616_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10003_ (.A1(_01940_),
    .A2(_04615_),
    .B(_04617_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10004_ (.A1(\as2650.stack[4][13] ),
    .A2(_04616_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10005_ (.A1(_01947_),
    .A2(_04615_),
    .B(_04618_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10006_ (.A1(\as2650.stack[4][14] ),
    .A2(_04616_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10007_ (.A1(_01954_),
    .A2(_04615_),
    .B(_04619_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10008_ (.A1(\as2650.stack[4][15] ),
    .A2(_04616_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10009_ (.A1(_01959_),
    .A2(_04615_),
    .B(_04620_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10010_ (.I(_01736_),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10011_ (.I(_02537_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10012_ (.A1(_01961_),
    .A2(_01962_),
    .A3(_04622_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10013_ (.I(_04623_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10014_ (.I(_04624_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10015_ (.I(_04623_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10016_ (.I(_04626_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10017_ (.A1(\as2650.stack[10][0] ),
    .A2(_04627_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10018_ (.A1(_04621_),
    .A2(_04625_),
    .B(_04628_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10019_ (.I(_01759_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10020_ (.A1(\as2650.stack[10][1] ),
    .A2(_04627_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10021_ (.A1(_04629_),
    .A2(_04625_),
    .B(_04630_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10022_ (.I(_01776_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10023_ (.A1(\as2650.stack[10][2] ),
    .A2(_04627_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10024_ (.A1(_04631_),
    .A2(_04625_),
    .B(_04632_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10025_ (.I(_01800_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10026_ (.A1(\as2650.stack[10][3] ),
    .A2(_04627_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10027_ (.A1(_04633_),
    .A2(_04625_),
    .B(_04634_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10028_ (.I(_01819_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10029_ (.I(_04624_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10030_ (.I(_04626_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10031_ (.A1(\as2650.stack[10][4] ),
    .A2(_04637_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10032_ (.A1(_04635_),
    .A2(_04636_),
    .B(_04638_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10033_ (.I(_01834_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10034_ (.A1(\as2650.stack[10][5] ),
    .A2(_04637_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10035_ (.A1(_04639_),
    .A2(_04636_),
    .B(_04640_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10036_ (.I(_01852_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10037_ (.A1(\as2650.stack[10][6] ),
    .A2(_04637_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10038_ (.A1(_04641_),
    .A2(_04636_),
    .B(_04642_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10039_ (.I(_01868_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10040_ (.A1(\as2650.stack[10][7] ),
    .A2(_04637_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10041_ (.A1(_04643_),
    .A2(_04636_),
    .B(_04644_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10042_ (.I(_01882_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10043_ (.I(_04624_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10044_ (.I(_04626_),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10045_ (.A1(\as2650.stack[10][8] ),
    .A2(_04647_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10046_ (.A1(_04645_),
    .A2(_04646_),
    .B(_04648_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10047_ (.I(_01898_),
    .Z(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10048_ (.A1(\as2650.stack[10][9] ),
    .A2(_04647_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10049_ (.A1(_04649_),
    .A2(_04646_),
    .B(_04650_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10050_ (.I(_01912_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10051_ (.A1(\as2650.stack[10][10] ),
    .A2(_04647_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10052_ (.A1(_04651_),
    .A2(_04646_),
    .B(_04652_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10053_ (.I(_01927_),
    .Z(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10054_ (.A1(\as2650.stack[10][11] ),
    .A2(_04647_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10055_ (.A1(_04653_),
    .A2(_04646_),
    .B(_04654_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10056_ (.I(_01939_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10057_ (.I(_04624_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10058_ (.I(_04626_),
    .Z(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10059_ (.A1(\as2650.stack[10][12] ),
    .A2(_04657_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10060_ (.A1(_04655_),
    .A2(_04656_),
    .B(_04658_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10061_ (.I(_01946_),
    .Z(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10062_ (.A1(\as2650.stack[10][13] ),
    .A2(_04657_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10063_ (.A1(_04659_),
    .A2(_04656_),
    .B(_04660_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10064_ (.I(_01953_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10065_ (.A1(\as2650.stack[10][14] ),
    .A2(_04657_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10066_ (.A1(_04661_),
    .A2(_04656_),
    .B(_04662_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10067_ (.I(_01958_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10068_ (.A1(\as2650.stack[10][15] ),
    .A2(_04657_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10069_ (.A1(_04663_),
    .A2(_04656_),
    .B(_04664_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10070_ (.I(_02545_),
    .Z(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10071_ (.A1(_01961_),
    .A2(_01970_),
    .A3(_04665_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10072_ (.I(_04666_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10073_ (.I(_04667_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10074_ (.I(_04666_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10075_ (.I(_04669_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10076_ (.A1(\as2650.stack[3][0] ),
    .A2(_04670_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10077_ (.A1(_04621_),
    .A2(_04668_),
    .B(_04671_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10078_ (.A1(\as2650.stack[3][1] ),
    .A2(_04670_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10079_ (.A1(_04629_),
    .A2(_04668_),
    .B(_04672_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10080_ (.A1(\as2650.stack[3][2] ),
    .A2(_04670_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10081_ (.A1(_04631_),
    .A2(_04668_),
    .B(_04673_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10082_ (.A1(\as2650.stack[3][3] ),
    .A2(_04670_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10083_ (.A1(_04633_),
    .A2(_04668_),
    .B(_04674_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10084_ (.I(_04667_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10085_ (.I(_04669_),
    .Z(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10086_ (.A1(\as2650.stack[3][4] ),
    .A2(_04676_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10087_ (.A1(_04635_),
    .A2(_04675_),
    .B(_04677_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10088_ (.A1(\as2650.stack[3][5] ),
    .A2(_04676_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10089_ (.A1(_04639_),
    .A2(_04675_),
    .B(_04678_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10090_ (.A1(\as2650.stack[3][6] ),
    .A2(_04676_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10091_ (.A1(_04641_),
    .A2(_04675_),
    .B(_04679_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10092_ (.A1(\as2650.stack[3][7] ),
    .A2(_04676_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10093_ (.A1(_04643_),
    .A2(_04675_),
    .B(_04680_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10094_ (.I(_04667_),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10095_ (.I(_04669_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10096_ (.A1(\as2650.stack[3][8] ),
    .A2(_04682_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10097_ (.A1(_04645_),
    .A2(_04681_),
    .B(_04683_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10098_ (.A1(\as2650.stack[3][9] ),
    .A2(_04682_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10099_ (.A1(_04649_),
    .A2(_04681_),
    .B(_04684_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10100_ (.A1(\as2650.stack[3][10] ),
    .A2(_04682_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10101_ (.A1(_04651_),
    .A2(_04681_),
    .B(_04685_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10102_ (.A1(\as2650.stack[3][11] ),
    .A2(_04682_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10103_ (.A1(_04653_),
    .A2(_04681_),
    .B(_04686_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10104_ (.I(_04667_),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10105_ (.I(_04669_),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10106_ (.A1(\as2650.stack[3][12] ),
    .A2(_04688_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10107_ (.A1(_04655_),
    .A2(_04687_),
    .B(_04689_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10108_ (.A1(\as2650.stack[3][13] ),
    .A2(_04688_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10109_ (.A1(_04659_),
    .A2(_04687_),
    .B(_04690_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10110_ (.A1(\as2650.stack[3][14] ),
    .A2(_04688_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10111_ (.A1(_04661_),
    .A2(_04687_),
    .B(_04691_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10112_ (.A1(\as2650.stack[3][15] ),
    .A2(_04688_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10113_ (.A1(_04663_),
    .A2(_04687_),
    .B(_04692_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10114_ (.A1(_01228_),
    .A2(_03151_),
    .B(_04432_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10115_ (.A1(_01727_),
    .A2(_01697_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10116_ (.A1(_04693_),
    .A2(_04694_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10117_ (.A1(_01292_),
    .A2(_01243_),
    .A3(_03715_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10118_ (.A1(_01083_),
    .A2(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10119_ (.A1(_01606_),
    .A2(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10120_ (.A1(_03159_),
    .A2(_04698_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10121_ (.A1(_03812_),
    .A2(_04699_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10122_ (.I(_01502_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10123_ (.A1(_02714_),
    .A2(_01279_),
    .A3(_01508_),
    .A4(_02581_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10124_ (.I(_04702_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10125_ (.A1(_04701_),
    .A2(_04703_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10126_ (.A1(_01478_),
    .A2(_01503_),
    .A3(_03715_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10127_ (.A1(_01695_),
    .A2(_04373_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10128_ (.A1(\as2650.cycle[10] ),
    .A2(_01695_),
    .A3(_01528_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10129_ (.A1(_04704_),
    .A2(_04705_),
    .A3(_04706_),
    .A4(_04707_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10130_ (.A1(_01083_),
    .A2(_01573_),
    .A3(_03742_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _10131_ (.A1(_01262_),
    .A2(_01297_),
    .A3(_01318_),
    .A4(_01471_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10132_ (.A1(_01461_),
    .A2(_04701_),
    .A3(_04710_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10133_ (.A1(_01461_),
    .A2(_01483_),
    .A3(_04701_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10134_ (.A1(_04711_),
    .A2(_04712_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10135_ (.A1(_04697_),
    .A2(_04708_),
    .A3(_04709_),
    .A4(_04713_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10136_ (.A1(_01208_),
    .A2(_04185_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10137_ (.A1(_01182_),
    .A2(_01169_),
    .B1(_01425_),
    .B2(_01442_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10138_ (.A1(_04716_),
    .A2(_04715_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10139_ (.A1(_01082_),
    .A2(_01573_),
    .A3(_03743_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10140_ (.A1(_01695_),
    .A2(_02917_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10141_ (.A1(_01728_),
    .A2(_04717_),
    .B(_04718_),
    .C(_04719_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10142_ (.A1(_04714_),
    .A2(_04720_),
    .B(_02580_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10143_ (.A1(_04698_),
    .A2(_04721_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10144_ (.A1(_04695_),
    .A2(_04700_),
    .A3(_04722_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10145_ (.I(_04723_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10146_ (.A1(_04234_),
    .A2(_04236_),
    .A3(_04237_),
    .A4(_04238_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10147_ (.I(_04697_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10148_ (.I(_04706_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10149_ (.I(_04727_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10150_ (.I(_04705_),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10151_ (.A1(_01237_),
    .A2(_01099_),
    .A3(_03727_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10152_ (.I(_04730_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10153_ (.A1(_01082_),
    .A2(_01572_),
    .A3(_04715_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10154_ (.I(_04732_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10155_ (.I(_04702_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10156_ (.A1(_01411_),
    .A2(_01504_),
    .A3(_04734_),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10157_ (.I(_01503_),
    .Z(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10158_ (.I(_04703_),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10159_ (.A1(_04736_),
    .A2(_04737_),
    .B(_01412_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10160_ (.A1(_01237_),
    .A2(_01099_),
    .A3(_04186_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10161_ (.I(_04739_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10162_ (.A1(_04733_),
    .A2(_04735_),
    .A3(_04738_),
    .B1(_04740_),
    .B2(_03658_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10163_ (.I(_04730_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10164_ (.A1(_01615_),
    .A2(_04742_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10165_ (.I(_04718_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10166_ (.A1(_04731_),
    .A2(_04741_),
    .B(_04743_),
    .C(_04744_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10167_ (.I(_04705_),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10168_ (.A1(_04287_),
    .A2(_04744_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10169_ (.A1(_04746_),
    .A2(_04747_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _10170_ (.A1(_04239_),
    .A2(_04729_),
    .B1(_04745_),
    .B2(_04748_),
    .C(_04711_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10171_ (.I(_04719_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10172_ (.A1(_01412_),
    .A2(_04711_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10173_ (.A1(_04750_),
    .A2(_04751_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10174_ (.A1(_02893_),
    .A2(\as2650.instruction_args_latch[14] ),
    .B(_02474_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10175_ (.A1(_02922_),
    .A2(_04753_),
    .Z(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10176_ (.A1(_03741_),
    .A2(_04754_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10177_ (.I(_04719_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10178_ (.A1(_01165_),
    .A2(_02934_),
    .A3(_01795_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10179_ (.I(_04757_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10180_ (.A1(_04749_),
    .A2(_04752_),
    .B1(_04755_),
    .B2(_04756_),
    .C(_04758_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10181_ (.A1(_01412_),
    .A2(_04712_),
    .B(_04727_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10182_ (.I(_04707_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10183_ (.A1(_02659_),
    .A2(_04728_),
    .B1(_04759_),
    .B2(_04760_),
    .C(_04761_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10184_ (.I(_04697_),
    .Z(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10185_ (.I(_04707_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10186_ (.A1(_04387_),
    .A2(_04764_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10187_ (.A1(_04763_),
    .A2(_04765_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10188_ (.A1(_04725_),
    .A2(_04726_),
    .B1(_04762_),
    .B2(_04766_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10189_ (.I(_04767_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10190_ (.I(_03816_),
    .Z(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10191_ (.A1(_04769_),
    .A2(_04695_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10192_ (.I(_04770_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10193_ (.A1(_01727_),
    .A2(_01750_),
    .A3(_03735_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10194_ (.I(_04772_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10195_ (.I(_04773_),
    .Z(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10196_ (.I(_04773_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10197_ (.A1(_03475_),
    .A2(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10198_ (.A1(_01729_),
    .A2(_04188_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10199_ (.I(_04777_),
    .Z(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10200_ (.I(_04778_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10201_ (.A1(_03658_),
    .A2(_04774_),
    .B(_04776_),
    .C(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10202_ (.A1(_01697_),
    .A2(_04183_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10203_ (.I(_04781_),
    .Z(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10204_ (.I(_04782_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10205_ (.A1(_04167_),
    .A2(_04783_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10206_ (.A1(_04780_),
    .A2(_04784_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10207_ (.A1(_04700_),
    .A2(_04722_),
    .B(_04770_),
    .C(_04571_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10208_ (.I(_04786_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10209_ (.I(\as2650.regs[5][0] ),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10210_ (.A1(_04724_),
    .A2(_04768_),
    .B1(_04771_),
    .B2(_04785_),
    .C1(_04787_),
    .C2(_04788_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10211_ (.I(_04786_),
    .Z(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10212_ (.I(_01415_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10213_ (.I(_04757_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10214_ (.I(_04711_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10215_ (.I(_04744_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10216_ (.A1(_01194_),
    .A2(_02469_),
    .A3(_01696_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10217_ (.I(_04732_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10218_ (.I(_01503_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10219_ (.A1(_01372_),
    .A2(_04796_),
    .A3(_04737_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10220_ (.I(_04701_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10221_ (.I(_04703_),
    .Z(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10222_ (.A1(_04798_),
    .A2(_04799_),
    .B(_01415_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10223_ (.I(_04739_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10224_ (.A1(_04795_),
    .A2(_04797_),
    .A3(_04800_),
    .B1(_04801_),
    .B2(_01747_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10225_ (.A1(_01237_),
    .A2(_01099_),
    .A3(_01182_),
    .A4(_01169_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10226_ (.A1(_01568_),
    .A2(_01614_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10227_ (.A1(_04803_),
    .A2(_04804_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10228_ (.I(_04730_),
    .Z(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10229_ (.A1(_04794_),
    .A2(_04802_),
    .B(_04805_),
    .C(_04806_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10230_ (.I(_04709_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10231_ (.A1(_04358_),
    .A2(_04808_),
    .B(_04793_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10232_ (.A1(_01460_),
    .A2(_01795_),
    .A3(_02585_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10233_ (.I(_04810_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10234_ (.A1(_01599_),
    .A2(_04793_),
    .B1(_04807_),
    .B2(_04809_),
    .C(_04811_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10235_ (.A1(_04247_),
    .A2(_04729_),
    .B(_04792_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10236_ (.A1(_01238_),
    .A2(_02917_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10237_ (.I(_04814_),
    .Z(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10238_ (.A1(_01415_),
    .A2(_04792_),
    .B1(_04812_),
    .B2(_04813_),
    .C(_04815_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10239_ (.A1(_02922_),
    .A2(_04753_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10240_ (.I(_04817_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10241_ (.I(_04817_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10242_ (.A1(_02913_),
    .A2(_02927_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10243_ (.A1(_01413_),
    .A2(_04820_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10244_ (.A1(_04819_),
    .A2(_04821_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10245_ (.A1(_01616_),
    .A2(_04818_),
    .B(_04822_),
    .C(_04815_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10246_ (.A1(_04791_),
    .A2(_04823_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10247_ (.A1(_01083_),
    .A2(_04372_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10248_ (.I(_04825_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10249_ (.A1(_04790_),
    .A2(_04791_),
    .B1(_04816_),
    .B2(_04824_),
    .C(_04826_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10250_ (.A1(_02677_),
    .A2(_04728_),
    .B(_04761_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10251_ (.A1(_04382_),
    .A2(_04761_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10252_ (.A1(_01084_),
    .A2(_04696_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10253_ (.I(_04830_),
    .Z(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10254_ (.A1(_04827_),
    .A2(_04828_),
    .B(_04829_),
    .C(_04831_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10255_ (.A1(_04247_),
    .A2(_04831_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10256_ (.A1(_04832_),
    .A2(_04833_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10257_ (.I(_04723_),
    .Z(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10258_ (.A1(_03498_),
    .A2(_04775_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10259_ (.A1(_01747_),
    .A2(_04774_),
    .B(_04836_),
    .C(_04779_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10260_ (.A1(_04166_),
    .A2(_04783_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10261_ (.A1(_04837_),
    .A2(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10262_ (.I(_04770_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10263_ (.A1(_00863_),
    .A2(_04789_),
    .B1(_04834_),
    .B2(_04835_),
    .C1(_04839_),
    .C2(_04840_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10264_ (.I(\as2650.regs[5][2] ),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10265_ (.I(_04231_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10266_ (.I(_04763_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10267_ (.I(_04763_),
    .Z(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10268_ (.A1(_01084_),
    .A2(_04380_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10269_ (.I(_04845_),
    .Z(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10270_ (.A1(_01728_),
    .A2(_03730_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10271_ (.I(_04847_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10272_ (.I(_04803_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10273_ (.A1(_04736_),
    .A2(_04737_),
    .B(_01410_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10274_ (.A1(_04358_),
    .A2(_04796_),
    .A3(_04734_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10275_ (.A1(_04733_),
    .A2(_04850_),
    .A3(_04851_),
    .B1(_04740_),
    .B2(_01769_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10276_ (.I(_04803_),
    .Z(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10277_ (.A1(\as2650.debug_psl[5] ),
    .A2(_01614_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10278_ (.A1(_01625_),
    .A2(_04854_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10279_ (.A1(_04853_),
    .A2(_04855_),
    .B(_04742_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10280_ (.A1(_04849_),
    .A2(_04852_),
    .B(_04856_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10281_ (.I(_04847_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10282_ (.A1(_04360_),
    .A2(_04806_),
    .B(_04858_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10283_ (.A1(_01616_),
    .A2(_04848_),
    .B1(_04857_),
    .B2(_04859_),
    .C(_04746_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10284_ (.I(_04810_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10285_ (.A1(_04231_),
    .A2(_04861_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10286_ (.A1(_04860_),
    .A2(_04862_),
    .B(_04756_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10287_ (.I(_04754_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10288_ (.A1(_02893_),
    .A2(_02905_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10289_ (.A1(_02894_),
    .A2(_01406_),
    .B1(_01408_),
    .B2(_04865_),
    .C(_04754_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10290_ (.A1(_01626_),
    .A2(_04864_),
    .B(_04866_),
    .C(_04719_),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10291_ (.A1(_04712_),
    .A2(_04867_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10292_ (.A1(_01410_),
    .A2(_04758_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10293_ (.A1(_04863_),
    .A2(_04868_),
    .B(_04869_),
    .C(_04727_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10294_ (.A1(_02716_),
    .A2(_04826_),
    .B(_04845_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10295_ (.A1(_04385_),
    .A2(_04846_),
    .B1(_04870_),
    .B2(_04871_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10296_ (.A1(_04844_),
    .A2(_04872_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10297_ (.A1(_04842_),
    .A2(_04843_),
    .B(_04873_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10298_ (.A1(_03528_),
    .A2(_04775_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10299_ (.I(_04778_),
    .Z(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10300_ (.A1(_01769_),
    .A2(_04774_),
    .B(_04875_),
    .C(_04876_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10301_ (.A1(_04164_),
    .A2(_04783_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10302_ (.A1(_04877_),
    .A2(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10303_ (.A1(_04841_),
    .A2(_04789_),
    .B1(_04874_),
    .B2(_04835_),
    .C1(_04879_),
    .C2(_04840_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10304_ (.I(\as2650.regs[5][3] ),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10305_ (.I(_04224_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10306_ (.I(_04757_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10307_ (.I(_04703_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10308_ (.A1(_04736_),
    .A2(_04883_),
    .B(_01404_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10309_ (.A1(_01401_),
    .A2(_01504_),
    .A3(_04734_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10310_ (.A1(_04733_),
    .A2(_04884_),
    .A3(_04885_),
    .B1(_04740_),
    .B2(_04194_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10311_ (.A1(_04358_),
    .A2(_01372_),
    .B(\as2650.debug_psl[5] ),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10312_ (.A1(_01637_),
    .A2(_04887_),
    .Z(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10313_ (.A1(_04853_),
    .A2(_04888_),
    .B(_04742_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10314_ (.A1(_04849_),
    .A2(_04886_),
    .B(_04889_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10315_ (.A1(_03858_),
    .A2(_04806_),
    .B(_04858_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10316_ (.A1(_01626_),
    .A2(_04848_),
    .B1(_04890_),
    .B2(_04891_),
    .C(_04746_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10317_ (.A1(_04224_),
    .A2(_04861_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10318_ (.A1(_04892_),
    .A2(_04893_),
    .B(_04750_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10319_ (.A1(_02894_),
    .A2(_01402_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10320_ (.A1(_01399_),
    .A2(_04820_),
    .B(_04895_),
    .C(_04819_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10321_ (.A1(_04360_),
    .A2(_04818_),
    .B(_04896_),
    .C(_04814_),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10322_ (.I(_04825_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10323_ (.A1(_01404_),
    .A2(_04758_),
    .B(_04898_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10324_ (.A1(_04882_),
    .A2(_04894_),
    .A3(_04897_),
    .B(_04899_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10325_ (.A1(_02731_),
    .A2(_04898_),
    .B(_04845_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10326_ (.A1(_04390_),
    .A2(_04846_),
    .B1(_04900_),
    .B2(_04901_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10327_ (.A1(_04844_),
    .A2(_04902_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10328_ (.A1(_04881_),
    .A2(_04843_),
    .B(_04903_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10329_ (.A1(_03548_),
    .A2(_04775_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10330_ (.A1(_04194_),
    .A2(_04774_),
    .B(_04905_),
    .C(_04876_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10331_ (.A1(_04160_),
    .A2(_04783_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10332_ (.A1(_04906_),
    .A2(_04907_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10333_ (.A1(_04880_),
    .A2(_04789_),
    .B1(_04904_),
    .B2(_04835_),
    .C1(_04908_),
    .C2(_04840_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10334_ (.I(\as2650.regs[5][4] ),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10335_ (.I(_03847_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10336_ (.A1(_01389_),
    .A2(_04798_),
    .A3(_04799_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10337_ (.A1(_01505_),
    .A2(_04799_),
    .B(_01397_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10338_ (.A1(_04795_),
    .A2(_04911_),
    .A3(_04912_),
    .B1(_04801_),
    .B2(_00923_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10339_ (.A1(_01656_),
    .A2(_04808_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10340_ (.A1(_04808_),
    .A2(_04913_),
    .B(_04914_),
    .C(_04848_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10341_ (.A1(_04360_),
    .A2(_04793_),
    .B(_04811_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _10342_ (.A1(_01461_),
    .A2(_01505_),
    .A3(_04710_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10343_ (.A1(_04910_),
    .A2(_04861_),
    .B1(_04915_),
    .B2(_04916_),
    .C(_04917_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10344_ (.A1(_01397_),
    .A2(_04917_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10345_ (.A1(_04815_),
    .A2(_04919_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10346_ (.A1(_02894_),
    .A2(_01393_),
    .B1(_04865_),
    .B2(_01395_),
    .C(_04864_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10347_ (.A1(_03858_),
    .A2(_04819_),
    .B(_04814_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10348_ (.A1(_04921_),
    .A2(_04922_),
    .B(_04882_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10349_ (.A1(_04918_),
    .A2(_04920_),
    .B(_04923_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10350_ (.A1(_01397_),
    .A2(_04791_),
    .B(_04826_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10351_ (.A1(_02626_),
    .A2(_04728_),
    .B(_04764_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10352_ (.A1(_04924_),
    .A2(_04925_),
    .B(_04926_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10353_ (.A1(_04386_),
    .A2(_04846_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10354_ (.A1(_04927_),
    .A2(_04928_),
    .B(_04831_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10355_ (.A1(_03847_),
    .A2(_04844_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10356_ (.A1(_04929_),
    .A2(_04930_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10357_ (.I(_04773_),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10358_ (.I(_04772_),
    .Z(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10359_ (.I(_04933_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10360_ (.A1(_03573_),
    .A2(_04934_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10361_ (.A1(_01804_),
    .A2(_04932_),
    .B(_04935_),
    .C(_04876_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10362_ (.A1(_04162_),
    .A2(_04782_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10363_ (.A1(_04936_),
    .A2(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10364_ (.A1(_04909_),
    .A2(_04789_),
    .B1(_04931_),
    .B2(_04835_),
    .C1(_04938_),
    .C2(_04840_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10365_ (.I(\as2650.regs[5][5] ),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10366_ (.I(_01387_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10367_ (.A1(_04282_),
    .A2(_04796_),
    .A3(_04883_),
    .Z(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10368_ (.A1(_04798_),
    .A2(_04737_),
    .B(_01387_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10369_ (.A1(_04795_),
    .A2(_04941_),
    .A3(_04942_),
    .B1(_04801_),
    .B2(_01823_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10370_ (.A1(_01557_),
    .A2(_04282_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10371_ (.A1(_04803_),
    .A2(_04944_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10372_ (.A1(_04794_),
    .A2(_04943_),
    .B(_04945_),
    .C(_04731_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10373_ (.A1(_03856_),
    .A2(_04808_),
    .B(_04744_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10374_ (.A1(_01648_),
    .A2(_04793_),
    .B1(_04946_),
    .B2(_04947_),
    .C(_04811_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10375_ (.I(_04216_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10376_ (.A1(_04949_),
    .A2(_04729_),
    .B(_04792_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _10377_ (.A1(_01387_),
    .A2(_04792_),
    .B1(_04948_),
    .B2(_04950_),
    .C(_04815_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10378_ (.A1(_02893_),
    .A2(_01384_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10379_ (.A1(_01385_),
    .A2(_04820_),
    .B(_04952_),
    .C(_04817_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10380_ (.A1(_01657_),
    .A2(_04818_),
    .B(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10381_ (.A1(_04756_),
    .A2(_04954_),
    .B(_04882_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10382_ (.A1(_04940_),
    .A2(_04791_),
    .B1(_04951_),
    .B2(_04955_),
    .C(_04826_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10383_ (.A1(_02781_),
    .A2(_04728_),
    .B(_04761_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10384_ (.A1(_04388_),
    .A2(_04764_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10385_ (.A1(_04956_),
    .A2(_04957_),
    .B(_04958_),
    .C(_04831_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10386_ (.A1(_04216_),
    .A2(_04726_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10387_ (.A1(_04959_),
    .A2(_04960_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10388_ (.A1(_02553_),
    .A2(_04934_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10389_ (.I(_04777_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10390_ (.I(_04963_),
    .Z(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10391_ (.A1(_01823_),
    .A2(_04932_),
    .B(_04962_),
    .C(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10392_ (.A1(_04159_),
    .A2(_04779_),
    .B(_04965_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10393_ (.A1(_04939_),
    .A2(_04787_),
    .B1(_04961_),
    .B2(_04724_),
    .C1(_04966_),
    .C2(_04771_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10394_ (.I(\as2650.regs[5][6] ),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10395_ (.A1(_04736_),
    .A2(_04883_),
    .B(_01423_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10396_ (.A1(_03856_),
    .A2(_01504_),
    .A3(_04734_),
    .Z(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10397_ (.A1(_04733_),
    .A2(_04968_),
    .A3(_04969_),
    .B1(_04740_),
    .B2(_01837_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10398_ (.A1(_01557_),
    .A2(_01383_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10399_ (.A1(_03855_),
    .A2(_04971_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10400_ (.A1(_04853_),
    .A2(_04972_),
    .B(_04742_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10401_ (.A1(_04849_),
    .A2(_04970_),
    .B(_04973_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10402_ (.A1(_03745_),
    .A2(_04731_),
    .B(_04847_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10403_ (.A1(_01657_),
    .A2(_04858_),
    .B1(_04974_),
    .B2(_04975_),
    .C(_04746_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10404_ (.A1(_04210_),
    .A2(_04811_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10405_ (.A1(_04976_),
    .A2(_04977_),
    .B(_04750_),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10406_ (.A1(_03036_),
    .A2(_01421_),
    .B1(_01420_),
    .B2(_04820_),
    .C(_04819_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10407_ (.A1(_03857_),
    .A2(_04818_),
    .B(_04979_),
    .C(_04814_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10408_ (.A1(_01423_),
    .A2(_04758_),
    .B(_04898_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10409_ (.A1(_04882_),
    .A2(_04978_),
    .A3(_04980_),
    .B(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10410_ (.A1(_02790_),
    .A2(_04898_),
    .B(_04845_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10411_ (.A1(_04389_),
    .A2(_04846_),
    .B1(_04982_),
    .B2(_04983_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10412_ (.A1(_04726_),
    .A2(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10413_ (.A1(_04364_),
    .A2(_04843_),
    .B(_04985_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10414_ (.A1(_03120_),
    .A2(_04934_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10415_ (.A1(_01838_),
    .A2(_04932_),
    .B(_04987_),
    .C(_04964_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10416_ (.A1(_04157_),
    .A2(_04779_),
    .B(_04988_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10417_ (.A1(_04967_),
    .A2(_04787_),
    .B1(_04986_),
    .B2(_04724_),
    .C1(_04989_),
    .C2(_04771_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10418_ (.I(\as2650.regs[5][7] ),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10419_ (.A1(_03744_),
    .A2(_04796_),
    .A3(_04883_),
    .Z(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10420_ (.A1(_04798_),
    .A2(_04799_),
    .B(_01382_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10421_ (.A1(_04795_),
    .A2(_04991_),
    .A3(_04992_),
    .B1(_04801_),
    .B2(_01856_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10422_ (.A1(_03855_),
    .A2(_01383_),
    .B(_03580_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10423_ (.A1(_00738_),
    .A2(_04994_),
    .Z(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10424_ (.A1(_04853_),
    .A2(_04995_),
    .B(_04731_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10425_ (.A1(_04849_),
    .A2(_04993_),
    .B(_04996_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10426_ (.A1(_04279_),
    .A2(_04806_),
    .B(_04858_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10427_ (.A1(_01664_),
    .A2(_04848_),
    .B1(_04997_),
    .B2(_04998_),
    .C(_04729_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10428_ (.A1(_03783_),
    .A2(_04861_),
    .B(_04917_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10429_ (.A1(_01382_),
    .A2(_04917_),
    .B1(_04999_),
    .B2(_05000_),
    .C(_04756_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10430_ (.A1(_02913_),
    .A2(_01363_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10431_ (.A1(_01380_),
    .A2(_04865_),
    .B(_05002_),
    .C(_04864_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10432_ (.A1(_01674_),
    .A2(_04864_),
    .B(_05003_),
    .C(_04750_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10433_ (.A1(_04727_),
    .A2(_05004_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10434_ (.A1(_01085_),
    .A2(_04426_),
    .B1(_05001_),
    .B2(_05005_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10435_ (.A1(_04393_),
    .A2(_04764_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10436_ (.A1(_04763_),
    .A2(_05007_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10437_ (.A1(_04365_),
    .A2(_04830_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10438_ (.A1(_05006_),
    .A2(_05008_),
    .B(_05009_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10439_ (.I(_05010_),
    .Z(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10440_ (.A1(_03146_),
    .A2(_04934_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10441_ (.A1(_01857_),
    .A2(_04932_),
    .B(_05012_),
    .C(_04876_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10442_ (.A1(_04156_),
    .A2(_04782_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10443_ (.A1(_05013_),
    .A2(_05014_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10444_ (.A1(_04990_),
    .A2(_04787_),
    .B1(_05011_),
    .B2(_04724_),
    .C1(_05015_),
    .C2(_04771_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10445_ (.I(_01712_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10446_ (.A1(_05016_),
    .A2(_04665_),
    .A3(_04622_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10447_ (.I(_05017_),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10448_ (.I(_05018_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10449_ (.I(_05017_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10450_ (.I(_05020_),
    .Z(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10451_ (.A1(\as2650.stack[2][0] ),
    .A2(_05021_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10452_ (.A1(_04621_),
    .A2(_05019_),
    .B(_05022_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10453_ (.A1(\as2650.stack[2][1] ),
    .A2(_05021_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10454_ (.A1(_04629_),
    .A2(_05019_),
    .B(_05023_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10455_ (.A1(\as2650.stack[2][2] ),
    .A2(_05021_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10456_ (.A1(_04631_),
    .A2(_05019_),
    .B(_05024_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10457_ (.A1(\as2650.stack[2][3] ),
    .A2(_05021_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10458_ (.A1(_04633_),
    .A2(_05019_),
    .B(_05025_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10459_ (.I(_05018_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10460_ (.I(_05020_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10461_ (.A1(\as2650.stack[2][4] ),
    .A2(_05027_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10462_ (.A1(_04635_),
    .A2(_05026_),
    .B(_05028_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10463_ (.A1(\as2650.stack[2][5] ),
    .A2(_05027_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10464_ (.A1(_04639_),
    .A2(_05026_),
    .B(_05029_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10465_ (.A1(\as2650.stack[2][6] ),
    .A2(_05027_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10466_ (.A1(_04641_),
    .A2(_05026_),
    .B(_05030_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10467_ (.A1(\as2650.stack[2][7] ),
    .A2(_05027_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10468_ (.A1(_04643_),
    .A2(_05026_),
    .B(_05031_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10469_ (.I(_05018_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10470_ (.I(_05020_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10471_ (.A1(\as2650.stack[2][8] ),
    .A2(_05033_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10472_ (.A1(_04645_),
    .A2(_05032_),
    .B(_05034_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10473_ (.A1(\as2650.stack[2][9] ),
    .A2(_05033_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10474_ (.A1(_04649_),
    .A2(_05032_),
    .B(_05035_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10475_ (.A1(\as2650.stack[2][10] ),
    .A2(_05033_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10476_ (.A1(_04651_),
    .A2(_05032_),
    .B(_05036_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10477_ (.A1(\as2650.stack[2][11] ),
    .A2(_05033_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10478_ (.A1(_04653_),
    .A2(_05032_),
    .B(_05037_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10479_ (.I(_05018_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10480_ (.I(_05020_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10481_ (.A1(\as2650.stack[2][12] ),
    .A2(_05039_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10482_ (.A1(_04655_),
    .A2(_05038_),
    .B(_05040_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10483_ (.A1(\as2650.stack[2][13] ),
    .A2(_05039_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10484_ (.A1(_04659_),
    .A2(_05038_),
    .B(_05041_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10485_ (.A1(\as2650.stack[2][14] ),
    .A2(_05039_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10486_ (.A1(_04661_),
    .A2(_05038_),
    .B(_05042_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10487_ (.A1(\as2650.stack[2][15] ),
    .A2(_05039_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10488_ (.A1(_04663_),
    .A2(_05038_),
    .B(_05043_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10489_ (.A1(_05016_),
    .A2(_04665_),
    .A3(_04522_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10490_ (.I(_05044_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10491_ (.I(_05045_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10492_ (.I(_05044_),
    .Z(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10493_ (.I(_05047_),
    .Z(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10494_ (.A1(\as2650.stack[1][0] ),
    .A2(_05048_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10495_ (.A1(_04621_),
    .A2(_05046_),
    .B(_05049_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10496_ (.A1(\as2650.stack[1][1] ),
    .A2(_05048_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10497_ (.A1(_04629_),
    .A2(_05046_),
    .B(_05050_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10498_ (.A1(\as2650.stack[1][2] ),
    .A2(_05048_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10499_ (.A1(_04631_),
    .A2(_05046_),
    .B(_05051_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10500_ (.A1(\as2650.stack[1][3] ),
    .A2(_05048_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10501_ (.A1(_04633_),
    .A2(_05046_),
    .B(_05052_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10502_ (.I(_05045_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10503_ (.I(_05047_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10504_ (.A1(\as2650.stack[1][4] ),
    .A2(_05054_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10505_ (.A1(_04635_),
    .A2(_05053_),
    .B(_05055_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10506_ (.A1(\as2650.stack[1][5] ),
    .A2(_05054_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10507_ (.A1(_04639_),
    .A2(_05053_),
    .B(_05056_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10508_ (.A1(\as2650.stack[1][6] ),
    .A2(_05054_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10509_ (.A1(_04641_),
    .A2(_05053_),
    .B(_05057_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10510_ (.A1(\as2650.stack[1][7] ),
    .A2(_05054_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10511_ (.A1(_04643_),
    .A2(_05053_),
    .B(_05058_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10512_ (.I(_05045_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10513_ (.I(_05047_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10514_ (.A1(\as2650.stack[1][8] ),
    .A2(_05060_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10515_ (.A1(_04645_),
    .A2(_05059_),
    .B(_05061_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10516_ (.A1(\as2650.stack[1][9] ),
    .A2(_05060_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10517_ (.A1(_04649_),
    .A2(_05059_),
    .B(_05062_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10518_ (.A1(\as2650.stack[1][10] ),
    .A2(_05060_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10519_ (.A1(_04651_),
    .A2(_05059_),
    .B(_05063_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10520_ (.A1(\as2650.stack[1][11] ),
    .A2(_05060_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10521_ (.A1(_04653_),
    .A2(_05059_),
    .B(_05064_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10522_ (.I(_05045_),
    .Z(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10523_ (.I(_05047_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10524_ (.A1(\as2650.stack[1][12] ),
    .A2(_05066_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10525_ (.A1(_04655_),
    .A2(_05065_),
    .B(_05067_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10526_ (.A1(\as2650.stack[1][13] ),
    .A2(_05066_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10527_ (.A1(_04659_),
    .A2(_05065_),
    .B(_05068_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10528_ (.A1(\as2650.stack[1][14] ),
    .A2(_05066_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10529_ (.A1(_04661_),
    .A2(_05065_),
    .B(_05069_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10530_ (.A1(\as2650.stack[1][15] ),
    .A2(_05066_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10531_ (.A1(_04663_),
    .A2(_05065_),
    .B(_05070_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10532_ (.I(_01736_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10533_ (.A1(_01685_),
    .A2(_01713_),
    .A3(_01970_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10534_ (.I(_05072_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10535_ (.I(_05073_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10536_ (.I(_05072_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10537_ (.I(_05075_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10538_ (.A1(\as2650.stack[15][0] ),
    .A2(_05076_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10539_ (.A1(_05071_),
    .A2(_05074_),
    .B(_05077_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10540_ (.I(_01759_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10541_ (.A1(\as2650.stack[15][1] ),
    .A2(_05076_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10542_ (.A1(_05078_),
    .A2(_05074_),
    .B(_05079_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10543_ (.I(_01776_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10544_ (.A1(\as2650.stack[15][2] ),
    .A2(_05076_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10545_ (.A1(_05080_),
    .A2(_05074_),
    .B(_05081_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10546_ (.I(_01800_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10547_ (.A1(\as2650.stack[15][3] ),
    .A2(_05076_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10548_ (.A1(_05082_),
    .A2(_05074_),
    .B(_05083_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10549_ (.I(_01819_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10550_ (.I(_05073_),
    .Z(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10551_ (.I(_05075_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10552_ (.A1(\as2650.stack[15][4] ),
    .A2(_05086_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10553_ (.A1(_05084_),
    .A2(_05085_),
    .B(_05087_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10554_ (.I(_01834_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10555_ (.A1(\as2650.stack[15][5] ),
    .A2(_05086_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10556_ (.A1(_05088_),
    .A2(_05085_),
    .B(_05089_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10557_ (.I(_01852_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10558_ (.A1(\as2650.stack[15][6] ),
    .A2(_05086_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10559_ (.A1(_05090_),
    .A2(_05085_),
    .B(_05091_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10560_ (.I(_01868_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10561_ (.A1(\as2650.stack[15][7] ),
    .A2(_05086_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10562_ (.A1(_05092_),
    .A2(_05085_),
    .B(_05093_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10563_ (.I(_01882_),
    .Z(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10564_ (.I(_05073_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10565_ (.I(_05075_),
    .Z(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10566_ (.A1(\as2650.stack[15][8] ),
    .A2(_05096_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10567_ (.A1(_05094_),
    .A2(_05095_),
    .B(_05097_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10568_ (.I(_01898_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10569_ (.A1(\as2650.stack[15][9] ),
    .A2(_05096_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10570_ (.A1(_05098_),
    .A2(_05095_),
    .B(_05099_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10571_ (.I(_01912_),
    .Z(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10572_ (.A1(\as2650.stack[15][10] ),
    .A2(_05096_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10573_ (.A1(_05100_),
    .A2(_05095_),
    .B(_05101_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10574_ (.I(_01927_),
    .Z(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10575_ (.A1(\as2650.stack[15][11] ),
    .A2(_05096_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10576_ (.A1(_05102_),
    .A2(_05095_),
    .B(_05103_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10577_ (.I(_01939_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10578_ (.I(_05073_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10579_ (.I(_05075_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10580_ (.A1(\as2650.stack[15][12] ),
    .A2(_05106_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10581_ (.A1(_05104_),
    .A2(_05105_),
    .B(_05107_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10582_ (.I(_01946_),
    .Z(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10583_ (.A1(\as2650.stack[15][13] ),
    .A2(_05106_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10584_ (.A1(_05108_),
    .A2(_05105_),
    .B(_05109_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10585_ (.I(_01953_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10586_ (.A1(\as2650.stack[15][14] ),
    .A2(_05106_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10587_ (.A1(_05110_),
    .A2(_05105_),
    .B(_05111_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10588_ (.I(_01958_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10589_ (.A1(\as2650.stack[15][15] ),
    .A2(_05106_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10590_ (.A1(_05112_),
    .A2(_05105_),
    .B(_05113_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10591_ (.A1(_05016_),
    .A2(_01970_),
    .A3(_04523_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10592_ (.I(_05114_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10593_ (.I(_05115_),
    .Z(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10594_ (.I(_05114_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10595_ (.I(_05117_),
    .Z(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10596_ (.A1(\as2650.stack[7][0] ),
    .A2(_05118_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10597_ (.A1(_05071_),
    .A2(_05116_),
    .B(_05119_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10598_ (.A1(\as2650.stack[7][1] ),
    .A2(_05118_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10599_ (.A1(_05078_),
    .A2(_05116_),
    .B(_05120_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10600_ (.A1(\as2650.stack[7][2] ),
    .A2(_05118_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10601_ (.A1(_05080_),
    .A2(_05116_),
    .B(_05121_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10602_ (.A1(\as2650.stack[7][3] ),
    .A2(_05118_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10603_ (.A1(_05082_),
    .A2(_05116_),
    .B(_05122_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10604_ (.I(_05115_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10605_ (.I(_05117_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10606_ (.A1(\as2650.stack[7][4] ),
    .A2(_05124_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10607_ (.A1(_05084_),
    .A2(_05123_),
    .B(_05125_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10608_ (.A1(\as2650.stack[7][5] ),
    .A2(_05124_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10609_ (.A1(_05088_),
    .A2(_05123_),
    .B(_05126_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10610_ (.A1(\as2650.stack[7][6] ),
    .A2(_05124_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10611_ (.A1(_05090_),
    .A2(_05123_),
    .B(_05127_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10612_ (.A1(\as2650.stack[7][7] ),
    .A2(_05124_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10613_ (.A1(_05092_),
    .A2(_05123_),
    .B(_05128_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10614_ (.I(_05115_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10615_ (.I(_05117_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10616_ (.A1(\as2650.stack[7][8] ),
    .A2(_05130_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10617_ (.A1(_05094_),
    .A2(_05129_),
    .B(_05131_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10618_ (.A1(\as2650.stack[7][9] ),
    .A2(_05130_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10619_ (.A1(_05098_),
    .A2(_05129_),
    .B(_05132_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10620_ (.A1(\as2650.stack[7][10] ),
    .A2(_05130_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10621_ (.A1(_05100_),
    .A2(_05129_),
    .B(_05133_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10622_ (.A1(\as2650.stack[7][11] ),
    .A2(_05130_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10623_ (.A1(_05102_),
    .A2(_05129_),
    .B(_05134_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10624_ (.I(_05115_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10625_ (.I(_05117_),
    .Z(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10626_ (.A1(\as2650.stack[7][12] ),
    .A2(_05136_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10627_ (.A1(_05104_),
    .A2(_05135_),
    .B(_05137_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10628_ (.A1(\as2650.stack[7][13] ),
    .A2(_05136_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10629_ (.A1(_05108_),
    .A2(_05135_),
    .B(_05138_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10630_ (.A1(\as2650.stack[7][14] ),
    .A2(_05136_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10631_ (.A1(_05110_),
    .A2(_05135_),
    .B(_05139_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10632_ (.A1(\as2650.stack[7][15] ),
    .A2(_05136_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10633_ (.A1(_05112_),
    .A2(_05135_),
    .B(_05140_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10634_ (.I(_04698_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10635_ (.A1(_02590_),
    .A2(_05141_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10636_ (.A1(_01807_),
    .A2(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10637_ (.A1(_04698_),
    .A2(_04721_),
    .A3(_05143_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10638_ (.A1(_04695_),
    .A2(_05144_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10639_ (.I(_05145_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10640_ (.A1(_04693_),
    .A2(_04694_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10641_ (.A1(_01808_),
    .A2(_05147_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10642_ (.I(_05148_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10643_ (.A1(_04571_),
    .A2(_05144_),
    .A3(_05148_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10644_ (.I(_05150_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10645_ (.I(\as2650.regs[1][0] ),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _10646_ (.A1(_04768_),
    .A2(_05146_),
    .B1(_05149_),
    .B2(_04785_),
    .C1(_05151_),
    .C2(_05152_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10647_ (.I(\as2650.regs[1][1] ),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _10648_ (.A1(_04834_),
    .A2(_05146_),
    .B1(_05149_),
    .B2(_04839_),
    .C1(_05151_),
    .C2(_05153_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10649_ (.I(\as2650.regs[1][2] ),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10650_ (.A1(_04874_),
    .A2(_05146_),
    .B1(_05149_),
    .B2(_04879_),
    .C1(_05151_),
    .C2(_05154_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10651_ (.I(\as2650.regs[1][3] ),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10652_ (.A1(_04904_),
    .A2(_05146_),
    .B1(_05149_),
    .B2(_04908_),
    .C1(_05151_),
    .C2(_05155_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10653_ (.I(_05145_),
    .Z(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10654_ (.I(_05148_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10655_ (.I(_05150_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10656_ (.I(\as2650.regs[1][4] ),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10657_ (.A1(_04931_),
    .A2(_05156_),
    .B1(_05157_),
    .B2(_04938_),
    .C1(_05158_),
    .C2(_05159_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10658_ (.I(\as2650.regs[1][5] ),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10659_ (.A1(_04961_),
    .A2(_05156_),
    .B1(_05157_),
    .B2(_04966_),
    .C1(_05158_),
    .C2(_05160_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10660_ (.I(\as2650.regs[1][6] ),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10661_ (.A1(_04986_),
    .A2(_05156_),
    .B1(_05157_),
    .B2(_04989_),
    .C1(_05158_),
    .C2(_05161_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10662_ (.I(\as2650.regs[1][7] ),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _10663_ (.A1(_05011_),
    .A2(_05156_),
    .B1(_05157_),
    .B2(_05015_),
    .C1(_05158_),
    .C2(_05162_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10664_ (.I(_04768_),
    .Z(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10665_ (.A1(_04714_),
    .A2(_04720_),
    .B(_04307_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10666_ (.A1(_01808_),
    .A2(_04699_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10667_ (.A1(_05164_),
    .A2(_05165_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10668_ (.I(_05166_),
    .Z(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10669_ (.I(_01240_),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10670_ (.A1(_05168_),
    .A2(_05166_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10671_ (.I(_05169_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10672_ (.A1(_05163_),
    .A2(_05167_),
    .B1(_05170_),
    .B2(_00848_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10673_ (.I(_04834_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10674_ (.A1(_05171_),
    .A2(_05167_),
    .B1(_05170_),
    .B2(_00867_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10675_ (.I(_04874_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10676_ (.A1(_05172_),
    .A2(_05167_),
    .B1(_05170_),
    .B2(_00890_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10677_ (.I(_04904_),
    .Z(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10678_ (.A1(_05173_),
    .A2(_05167_),
    .B1(_05170_),
    .B2(_00818_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10679_ (.I(_04931_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10680_ (.I(_05166_),
    .Z(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10681_ (.I(_05169_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10682_ (.A1(_05174_),
    .A2(_05175_),
    .B1(_05176_),
    .B2(_00916_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10683_ (.I(_04961_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10684_ (.A1(_05177_),
    .A2(_05175_),
    .B1(_05176_),
    .B2(_00795_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10685_ (.I(_04986_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10686_ (.A1(_05178_),
    .A2(_05175_),
    .B1(_05176_),
    .B2(_00759_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10687_ (.I(_05011_),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10688_ (.A1(_05179_),
    .A2(_05175_),
    .B1(_05176_),
    .B2(_00710_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10689_ (.A1(_04721_),
    .A2(_05165_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10690_ (.I(_05180_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10691_ (.A1(_05168_),
    .A2(_05180_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10692_ (.I(_05182_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10693_ (.A1(_05163_),
    .A2(_05181_),
    .B1(_05183_),
    .B2(_00842_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10694_ (.A1(_05171_),
    .A2(_05181_),
    .B1(_05183_),
    .B2(_00860_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10695_ (.A1(_05172_),
    .A2(_05181_),
    .B1(_05183_),
    .B2(_00884_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10696_ (.A1(_05173_),
    .A2(_05181_),
    .B1(_05183_),
    .B2(_00812_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10697_ (.I(_05180_),
    .Z(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10698_ (.I(_05182_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10699_ (.A1(_05174_),
    .A2(_05184_),
    .B1(_05185_),
    .B2(_00908_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10700_ (.A1(_05177_),
    .A2(_05184_),
    .B1(_05185_),
    .B2(_00785_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10701_ (.A1(_05178_),
    .A2(_05184_),
    .B1(_05185_),
    .B2(_00750_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10702_ (.A1(_05179_),
    .A2(_05184_),
    .B1(_05185_),
    .B2(_00695_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10703_ (.I(_01712_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10704_ (.A1(_01694_),
    .A2(_05186_),
    .A3(_01962_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10705_ (.I(_05187_),
    .Z(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10706_ (.I(_05188_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10707_ (.I(_05187_),
    .Z(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10708_ (.I(_05190_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10709_ (.A1(\as2650.stack[8][0] ),
    .A2(_05191_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10710_ (.A1(_05071_),
    .A2(_05189_),
    .B(_05192_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10711_ (.A1(\as2650.stack[8][1] ),
    .A2(_05191_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10712_ (.A1(_05078_),
    .A2(_05189_),
    .B(_05193_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10713_ (.A1(\as2650.stack[8][2] ),
    .A2(_05191_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10714_ (.A1(_05080_),
    .A2(_05189_),
    .B(_05194_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10715_ (.A1(\as2650.stack[8][3] ),
    .A2(_05191_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10716_ (.A1(_05082_),
    .A2(_05189_),
    .B(_05195_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10717_ (.I(_05188_),
    .Z(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10718_ (.I(_05190_),
    .Z(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10719_ (.A1(\as2650.stack[8][4] ),
    .A2(_05197_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10720_ (.A1(_05084_),
    .A2(_05196_),
    .B(_05198_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10721_ (.A1(\as2650.stack[8][5] ),
    .A2(_05197_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10722_ (.A1(_05088_),
    .A2(_05196_),
    .B(_05199_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10723_ (.A1(\as2650.stack[8][6] ),
    .A2(_05197_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10724_ (.A1(_05090_),
    .A2(_05196_),
    .B(_05200_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10725_ (.A1(\as2650.stack[8][7] ),
    .A2(_05197_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10726_ (.A1(_05092_),
    .A2(_05196_),
    .B(_05201_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10727_ (.I(_05188_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10728_ (.I(_05190_),
    .Z(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10729_ (.A1(\as2650.stack[8][8] ),
    .A2(_05203_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10730_ (.A1(_05094_),
    .A2(_05202_),
    .B(_05204_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10731_ (.A1(\as2650.stack[8][9] ),
    .A2(_05203_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10732_ (.A1(_05098_),
    .A2(_05202_),
    .B(_05205_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10733_ (.A1(\as2650.stack[8][10] ),
    .A2(_05203_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10734_ (.A1(_05100_),
    .A2(_05202_),
    .B(_05206_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(\as2650.stack[8][11] ),
    .A2(_05203_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10736_ (.A1(_05102_),
    .A2(_05202_),
    .B(_05207_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10737_ (.I(_05188_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10738_ (.I(_05190_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10739_ (.A1(\as2650.stack[8][12] ),
    .A2(_05209_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10740_ (.A1(_05104_),
    .A2(_05208_),
    .B(_05210_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10741_ (.A1(\as2650.stack[8][13] ),
    .A2(_05209_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10742_ (.A1(_05108_),
    .A2(_05208_),
    .B(_05211_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10743_ (.A1(\as2650.stack[8][14] ),
    .A2(_05209_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10744_ (.A1(_05110_),
    .A2(_05208_),
    .B(_05212_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10745_ (.A1(\as2650.stack[8][15] ),
    .A2(_05209_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10746_ (.A1(_05112_),
    .A2(_05208_),
    .B(_05213_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10747_ (.A1(_01584_),
    .A2(_01595_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10748_ (.A1(_04769_),
    .A2(_05142_),
    .A3(_05164_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10749_ (.I(_05214_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10750_ (.A1(_05168_),
    .A2(_05214_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10751_ (.I(_05216_),
    .Z(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10752_ (.I(\as2650.regs[6][0] ),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10753_ (.A1(_05163_),
    .A2(_05215_),
    .B1(_05217_),
    .B2(_05218_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10754_ (.I(\as2650.regs[6][1] ),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10755_ (.A1(_05171_),
    .A2(_05215_),
    .B1(_05217_),
    .B2(_05219_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10756_ (.I(\as2650.regs[6][2] ),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10757_ (.A1(_05172_),
    .A2(_05215_),
    .B1(_05217_),
    .B2(_05220_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10758_ (.I(\as2650.regs[6][3] ),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10759_ (.A1(_05173_),
    .A2(_05215_),
    .B1(_05217_),
    .B2(_05221_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10760_ (.I(_05214_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10761_ (.I(_05216_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10762_ (.I(\as2650.regs[6][4] ),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10763_ (.A1(_05174_),
    .A2(_05222_),
    .B1(_05223_),
    .B2(_05224_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10764_ (.I(\as2650.regs[6][5] ),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10765_ (.A1(_05177_),
    .A2(_05222_),
    .B1(_05223_),
    .B2(_05225_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10766_ (.I(\as2650.regs[6][6] ),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10767_ (.A1(_05178_),
    .A2(_05222_),
    .B1(_05223_),
    .B2(_05226_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10768_ (.I(\as2650.regs[6][7] ),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10769_ (.A1(_05179_),
    .A2(_05222_),
    .B1(_05223_),
    .B2(_05227_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10770_ (.A1(_05016_),
    .A2(_04622_),
    .A3(_04523_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10771_ (.I(_05228_),
    .Z(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10772_ (.I(_05229_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10773_ (.I(_05228_),
    .Z(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10774_ (.I(_05231_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10775_ (.A1(\as2650.stack[6][0] ),
    .A2(_05232_),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10776_ (.A1(_05071_),
    .A2(_05230_),
    .B(_05233_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10777_ (.A1(\as2650.stack[6][1] ),
    .A2(_05232_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10778_ (.A1(_05078_),
    .A2(_05230_),
    .B(_05234_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(\as2650.stack[6][2] ),
    .A2(_05232_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10780_ (.A1(_05080_),
    .A2(_05230_),
    .B(_05235_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10781_ (.A1(\as2650.stack[6][3] ),
    .A2(_05232_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10782_ (.A1(_05082_),
    .A2(_05230_),
    .B(_05236_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10783_ (.I(_05229_),
    .Z(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10784_ (.I(_05231_),
    .Z(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10785_ (.A1(\as2650.stack[6][4] ),
    .A2(_05238_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10786_ (.A1(_05084_),
    .A2(_05237_),
    .B(_05239_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10787_ (.A1(\as2650.stack[6][5] ),
    .A2(_05238_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10788_ (.A1(_05088_),
    .A2(_05237_),
    .B(_05240_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10789_ (.A1(\as2650.stack[6][6] ),
    .A2(_05238_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10790_ (.A1(_05090_),
    .A2(_05237_),
    .B(_05241_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10791_ (.A1(\as2650.stack[6][7] ),
    .A2(_05238_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10792_ (.A1(_05092_),
    .A2(_05237_),
    .B(_05242_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10793_ (.I(_05229_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10794_ (.I(_05231_),
    .Z(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10795_ (.A1(\as2650.stack[6][8] ),
    .A2(_05244_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10796_ (.A1(_05094_),
    .A2(_05243_),
    .B(_05245_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10797_ (.A1(\as2650.stack[6][9] ),
    .A2(_05244_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10798_ (.A1(_05098_),
    .A2(_05243_),
    .B(_05246_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10799_ (.A1(\as2650.stack[6][10] ),
    .A2(_05244_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10800_ (.A1(_05100_),
    .A2(_05243_),
    .B(_05247_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10801_ (.A1(\as2650.stack[6][11] ),
    .A2(_05244_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10802_ (.A1(_05102_),
    .A2(_05243_),
    .B(_05248_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10803_ (.I(_05229_),
    .Z(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10804_ (.I(_05231_),
    .Z(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10805_ (.A1(\as2650.stack[6][12] ),
    .A2(_05250_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10806_ (.A1(_05104_),
    .A2(_05249_),
    .B(_05251_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10807_ (.A1(\as2650.stack[6][13] ),
    .A2(_05250_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10808_ (.A1(_05108_),
    .A2(_05249_),
    .B(_05252_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10809_ (.A1(\as2650.stack[6][14] ),
    .A2(_05250_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10810_ (.A1(_05110_),
    .A2(_05249_),
    .B(_05253_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10811_ (.A1(\as2650.stack[6][15] ),
    .A2(_05250_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10812_ (.A1(_05112_),
    .A2(_05249_),
    .B(_05254_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10813_ (.A1(_01697_),
    .A2(_04300_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10814_ (.A1(_01579_),
    .A2(_01750_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10815_ (.A1(_01750_),
    .A2(_03725_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10816_ (.A1(_05255_),
    .A2(_05256_),
    .A3(_05257_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10817_ (.A1(_05147_),
    .A2(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10818_ (.A1(_03817_),
    .A2(_05259_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10819_ (.I(_05260_),
    .Z(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10820_ (.I(_05255_),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10821_ (.I(_05262_),
    .Z(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10822_ (.A1(_01492_),
    .A2(net219),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10823_ (.A1(_01749_),
    .A2(_01728_),
    .A3(_02476_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10824_ (.I(_05265_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10825_ (.I(_05256_),
    .Z(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10826_ (.A1(_03218_),
    .A2(_05266_),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10827_ (.A1(net219),
    .A2(_05266_),
    .B(_05267_),
    .C(_05268_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10828_ (.A1(_04187_),
    .A2(_01729_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10829_ (.I(_05270_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10830_ (.I(_04777_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10831_ (.A1(\as2650.chirpchar[0] ),
    .A2(_05271_),
    .B(_05272_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10832_ (.A1(_05264_),
    .A2(_04964_),
    .B1(_05269_),
    .B2(_05273_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10833_ (.I(_05257_),
    .Z(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10834_ (.I(_05275_),
    .Z(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10835_ (.I0(_05274_),
    .I1(_04725_),
    .S(_05276_),
    .Z(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10836_ (.A1(_03706_),
    .A2(_02580_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10837_ (.A1(_04440_),
    .A2(_02559_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10838_ (.I(_05262_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10839_ (.A1(_05278_),
    .A2(_05279_),
    .B(_05280_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10840_ (.A1(_05263_),
    .A2(_05277_),
    .B(_05281_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10841_ (.A1(_05141_),
    .A2(_05164_),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10842_ (.A1(_01807_),
    .A2(_04699_),
    .A3(_05283_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10843_ (.A1(_01085_),
    .A2(_05284_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10844_ (.A1(_05147_),
    .A2(_05258_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10845_ (.A1(_03812_),
    .A2(_05285_),
    .A3(_05286_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10846_ (.I(_05287_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10847_ (.A1(\as2650.regs[4][0] ),
    .A2(_05288_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10848_ (.I(_03812_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10849_ (.I(_05284_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10850_ (.A1(_05290_),
    .A2(_00851_),
    .A3(_01525_),
    .B1(_04767_),
    .B2(_05291_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10851_ (.A1(_05292_),
    .A2(_05260_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10852_ (.A1(_05261_),
    .A2(_05282_),
    .B(_05289_),
    .C(_05293_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10853_ (.A1(_03816_),
    .A2(_05259_),
    .Z(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10854_ (.I(_05294_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10855_ (.A1(_04832_),
    .A2(_04833_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10856_ (.I(_05284_),
    .Z(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10857_ (.I(_05285_),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10858_ (.A1(_05296_),
    .A2(_05297_),
    .B1(_05298_),
    .B2(_00871_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10859_ (.A1(\as2650.regs[4][1] ),
    .A2(_05288_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10860_ (.I(_05294_),
    .Z(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10861_ (.I(_05275_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10862_ (.I(_05275_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10863_ (.I(_05270_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10864_ (.A1(_01351_),
    .A2(_05265_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10865_ (.A1(_03268_),
    .A2(_05266_),
    .B(_05304_),
    .C(_05305_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10866_ (.A1(\as2650.chirpchar[1] ),
    .A2(_05267_),
    .B(_04781_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10867_ (.A1(_04038_),
    .A2(_04176_),
    .B(_04963_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10868_ (.A1(_05306_),
    .A2(_05307_),
    .B(_05308_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10869_ (.A1(_05303_),
    .A2(_05309_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10870_ (.A1(_04247_),
    .A2(_05302_),
    .B(_05310_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10871_ (.I(_05262_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10872_ (.I0(_05311_),
    .I1(_04318_),
    .S(_05312_),
    .Z(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10873_ (.A1(_05301_),
    .A2(_05313_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10874_ (.A1(_05295_),
    .A2(_05299_),
    .B(_05300_),
    .C(_05314_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10875_ (.I(_04726_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_04842_),
    .A2(_04844_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10877_ (.A1(_05315_),
    .A2(_04872_),
    .B(_05316_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10878_ (.A1(_05317_),
    .A2(_05284_),
    .B1(_05285_),
    .B2(_00894_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10879_ (.A1(\as2650.regs[4][2] ),
    .A2(_05288_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10880_ (.I(_05262_),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10881_ (.I(_05265_),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10882_ (.A1(_03311_),
    .A2(_05321_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10883_ (.A1(net189),
    .A2(_04933_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10884_ (.A1(_05322_),
    .A2(_05323_),
    .B(_05304_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10885_ (.A1(\as2650.chirpchar[2] ),
    .A2(_05271_),
    .B(_05324_),
    .C(_05272_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10886_ (.A1(_04175_),
    .A2(_04781_),
    .B(_05303_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10887_ (.A1(_04231_),
    .A2(_05276_),
    .B1(_05325_),
    .B2(_05326_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10888_ (.A1(_05320_),
    .A2(_05327_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10889_ (.A1(_04314_),
    .A2(_04315_),
    .A3(_05312_),
    .Z(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10890_ (.A1(_05328_),
    .A2(_05329_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10891_ (.A1(_05301_),
    .A2(_05330_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10892_ (.A1(_05301_),
    .A2(_05318_),
    .B(_05319_),
    .C(_05331_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10893_ (.A1(_04881_),
    .A2(_05315_),
    .ZN(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10894_ (.A1(_05315_),
    .A2(_04902_),
    .B(_05332_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10895_ (.A1(_05333_),
    .A2(_05297_),
    .B1(_05298_),
    .B2(_00822_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10896_ (.I(_05287_),
    .Z(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10897_ (.A1(_03335_),
    .A2(_05321_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10898_ (.A1(net190),
    .A2(_04933_),
    .B(_05304_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10899_ (.A1(\as2650.chirpchar[3] ),
    .A2(_05256_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10900_ (.A1(_05336_),
    .A2(_05337_),
    .B(_05338_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10901_ (.A1(_04174_),
    .A2(_04963_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10902_ (.I(_05275_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10903_ (.A1(_04778_),
    .A2(_05339_),
    .B(_05340_),
    .C(_05341_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10904_ (.A1(_04224_),
    .A2(_05302_),
    .B(_05342_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10905_ (.A1(_04310_),
    .A2(_05312_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10906_ (.A1(_05320_),
    .A2(_05343_),
    .B(_05344_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10907_ (.A1(_04480_),
    .A2(_02580_),
    .A3(_05280_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10908_ (.A1(_05345_),
    .A2(_05346_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10909_ (.A1(\as2650.regs[4][3] ),
    .A2(_05335_),
    .B1(_05347_),
    .B2(_05301_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10910_ (.A1(_05295_),
    .A2(_05334_),
    .B(_05348_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10911_ (.A1(_04929_),
    .A2(_04930_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10912_ (.A1(_05349_),
    .A2(_05297_),
    .B1(_05298_),
    .B2(_00921_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10913_ (.A1(_03362_),
    .A2(_05321_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10914_ (.A1(net191),
    .A2(_04772_),
    .B(_05270_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10915_ (.A1(\as2650.chirpchar[4] ),
    .A2(_05256_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10916_ (.A1(_05351_),
    .A2(_05352_),
    .B(_05353_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10917_ (.A1(_04173_),
    .A2(_04963_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10918_ (.A1(_05272_),
    .A2(_05354_),
    .B(_05355_),
    .C(_05341_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10919_ (.A1(_04910_),
    .A2(_05276_),
    .B(_05356_),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10920_ (.A1(_05320_),
    .A2(_05357_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10921_ (.A1(_04324_),
    .A2(_05263_),
    .B(_05358_),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10922_ (.A1(\as2650.regs[4][4] ),
    .A2(_05335_),
    .B1(_05359_),
    .B2(_05294_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10923_ (.A1(_05295_),
    .A2(_05350_),
    .B(_05360_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10924_ (.A1(_03386_),
    .A2(_05266_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10925_ (.A1(net192),
    .A2(_04933_),
    .B(_05271_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10926_ (.A1(\as2650.chirpchar[5] ),
    .A2(_05267_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10927_ (.A1(_05361_),
    .A2(_05362_),
    .B(_05363_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10928_ (.A1(_04171_),
    .A2(_04778_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10929_ (.A1(_04964_),
    .A2(_05364_),
    .B(_05365_),
    .C(_05276_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10930_ (.A1(_04949_),
    .A2(_05302_),
    .B(_05366_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10931_ (.A1(_04306_),
    .A2(_04308_),
    .A3(_05280_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10932_ (.A1(_05263_),
    .A2(_05367_),
    .B(_05368_),
    .ZN(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10933_ (.A1(\as2650.regs[4][5] ),
    .A2(_05288_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10934_ (.A1(_04959_),
    .A2(_04960_),
    .B(_05291_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10935_ (.A1(_05290_),
    .A2(_00801_),
    .A3(_01087_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10936_ (.A1(_05371_),
    .A2(_05372_),
    .B(_05260_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10937_ (.A1(_05261_),
    .A2(_05369_),
    .B(_05370_),
    .C(_05373_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10938_ (.A1(_04364_),
    .A2(_04843_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10939_ (.A1(_05315_),
    .A2(_04984_),
    .B(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10940_ (.A1(_05375_),
    .A2(_05297_),
    .B1(_05298_),
    .B2(_00763_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10941_ (.A1(_03416_),
    .A2(_05321_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10942_ (.A1(net193),
    .A2(_04772_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10943_ (.A1(_05377_),
    .A2(_05378_),
    .B(_05304_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10944_ (.A1(\as2650.chirpchar[6] ),
    .A2(_05271_),
    .B(_05379_),
    .C(_05272_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10945_ (.A1(_04169_),
    .A2(_04781_),
    .B(_05341_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10946_ (.A1(_04210_),
    .A2(_05303_),
    .B1(_05380_),
    .B2(_05381_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10947_ (.A1(_05320_),
    .A2(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10948_ (.A1(_04322_),
    .A2(_05280_),
    .B(_05383_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10949_ (.A1(\as2650.regs[4][6] ),
    .A2(_05335_),
    .B1(_05384_),
    .B2(_05294_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10950_ (.A1(_05295_),
    .A2(_05376_),
    .B(_05385_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10951_ (.A1(_03158_),
    .A2(_04432_),
    .A3(_03440_),
    .B(_04189_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10952_ (.A1(_01729_),
    .A2(_05386_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10953_ (.A1(net194),
    .A2(_04773_),
    .B(_05387_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10954_ (.A1(_04168_),
    .A2(_04782_),
    .B(_05303_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10955_ (.A1(_04365_),
    .A2(_05302_),
    .B1(_05388_),
    .B2(_05389_),
    .C(_05312_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10956_ (.A1(_04313_),
    .A2(_05263_),
    .B(_05390_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10957_ (.A1(\as2650.regs[4][7] ),
    .A2(_05335_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10958_ (.A1(_05290_),
    .A2(_00725_),
    .A3(_01525_),
    .B1(_05010_),
    .B2(_05291_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10959_ (.A1(_05261_),
    .A2(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10960_ (.A1(_05261_),
    .A2(_05391_),
    .B(_05392_),
    .C(_05394_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10961_ (.A1(_05255_),
    .A2(_05267_),
    .A3(_05341_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10962_ (.A1(_05147_),
    .A2(_05395_),
    .B(_03816_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10963_ (.I(_05396_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10964_ (.I(_05397_),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10965_ (.A1(_05143_),
    .A2(_05283_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10966_ (.A1(_03817_),
    .A2(\as2650.regs[4][0] ),
    .A3(_01547_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10967_ (.A1(_04768_),
    .A2(_05399_),
    .B(_05400_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10968_ (.A1(_05401_),
    .A2(_05398_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10969_ (.A1(_05143_),
    .A2(_05283_),
    .Z(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10970_ (.A1(_04769_),
    .A2(_01515_),
    .A3(_05259_),
    .A4(_05403_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10971_ (.I(_05404_),
    .Z(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10972_ (.A1(\as2650.regs[0][0] ),
    .A2(_05405_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10973_ (.A1(_05282_),
    .A2(_05398_),
    .B(_05402_),
    .C(_05406_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10974_ (.A1(_02201_),
    .A2(_05286_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10975_ (.I(_05407_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10976_ (.I(_05403_),
    .Z(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10977_ (.A1(_03813_),
    .A2(\as2650.regs[4][1] ),
    .A3(_03104_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10978_ (.A1(_05296_),
    .A2(_05409_),
    .B(_05410_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10979_ (.I(_05396_),
    .Z(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10980_ (.A1(_05313_),
    .A2(_05412_),
    .B1(_05405_),
    .B2(\as2650.regs[0][1] ),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10981_ (.A1(_05408_),
    .A2(_05411_),
    .B(_05413_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10982_ (.A1(_03813_),
    .A2(\as2650.regs[4][2] ),
    .A3(_03104_),
    .Z(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10983_ (.A1(_05317_),
    .A2(_05409_),
    .B(_05414_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10984_ (.I(_05404_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10985_ (.A1(_05330_),
    .A2(_05412_),
    .B1(_05416_),
    .B2(\as2650.regs[0][2] ),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10986_ (.A1(_05408_),
    .A2(_05415_),
    .B(_05417_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10987_ (.A1(_03813_),
    .A2(\as2650.regs[4][3] ),
    .A3(_02669_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10988_ (.A1(_05333_),
    .A2(_05409_),
    .B(_05418_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10989_ (.A1(_05347_),
    .A2(_05412_),
    .B1(_05416_),
    .B2(\as2650.regs[0][3] ),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10990_ (.A1(_05408_),
    .A2(_05419_),
    .B(_05420_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10991_ (.A1(_02201_),
    .A2(\as2650.regs[4][4] ),
    .A3(_02669_),
    .Z(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10992_ (.A1(_05349_),
    .A2(_05409_),
    .B(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10993_ (.A1(_05359_),
    .A2(_05412_),
    .B1(_05416_),
    .B2(\as2650.regs[0][4] ),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10994_ (.A1(_05408_),
    .A2(_05422_),
    .B(_05423_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10995_ (.A1(_04959_),
    .A2(_04960_),
    .B(_05399_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10996_ (.A1(_05290_),
    .A2(\as2650.regs[4][5] ),
    .A3(_03104_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10997_ (.A1(_05424_),
    .A2(_05425_),
    .B(_05397_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10998_ (.A1(\as2650.regs[0][5] ),
    .A2(_05405_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10999_ (.A1(_05369_),
    .A2(_05398_),
    .B(_05426_),
    .C(_05427_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11000_ (.A1(_03817_),
    .A2(\as2650.regs[4][6] ),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11001_ (.A1(_05428_),
    .A2(_01534_),
    .A3(_05403_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11002_ (.A1(_05375_),
    .A2(_05403_),
    .B(_05429_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11003_ (.A1(_05384_),
    .A2(_05396_),
    .B1(_05416_),
    .B2(\as2650.regs[0][6] ),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11004_ (.A1(_05407_),
    .A2(_05430_),
    .B(_05431_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11005_ (.A1(_02201_),
    .A2(\as2650.regs[4][7] ),
    .A3(_02669_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11006_ (.A1(_05011_),
    .A2(_05399_),
    .B(_05432_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11007_ (.A1(_05397_),
    .A2(_05433_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11008_ (.A1(\as2650.regs[0][7] ),
    .A2(_05405_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11009_ (.A1(_05391_),
    .A2(_05398_),
    .B(_05434_),
    .C(_05435_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11010_ (.I(_01736_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11011_ (.A1(_01694_),
    .A2(_05186_),
    .A3(_04665_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11012_ (.I(_05437_),
    .Z(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11013_ (.I(_05438_),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11014_ (.I(_05437_),
    .Z(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11015_ (.I(_05440_),
    .Z(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11016_ (.A1(\as2650.stack[0][0] ),
    .A2(_05441_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11017_ (.A1(_05436_),
    .A2(_05439_),
    .B(_05442_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11018_ (.I(_01759_),
    .Z(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11019_ (.A1(\as2650.stack[0][1] ),
    .A2(_05441_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11020_ (.A1(_05443_),
    .A2(_05439_),
    .B(_05444_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11021_ (.I(_01776_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11022_ (.A1(\as2650.stack[0][2] ),
    .A2(_05441_),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11023_ (.A1(_05445_),
    .A2(_05439_),
    .B(_05446_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11024_ (.I(_01800_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11025_ (.A1(\as2650.stack[0][3] ),
    .A2(_05441_),
    .ZN(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11026_ (.A1(_05447_),
    .A2(_05439_),
    .B(_05448_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11027_ (.I(_01819_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11028_ (.I(_05438_),
    .Z(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11029_ (.I(_05440_),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11030_ (.A1(\as2650.stack[0][4] ),
    .A2(_05451_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11031_ (.A1(_05449_),
    .A2(_05450_),
    .B(_05452_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11032_ (.I(_01834_),
    .Z(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11033_ (.A1(\as2650.stack[0][5] ),
    .A2(_05451_),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11034_ (.A1(_05453_),
    .A2(_05450_),
    .B(_05454_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11035_ (.I(_01852_),
    .Z(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11036_ (.A1(\as2650.stack[0][6] ),
    .A2(_05451_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11037_ (.A1(_05455_),
    .A2(_05450_),
    .B(_05456_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11038_ (.I(_01868_),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11039_ (.A1(\as2650.stack[0][7] ),
    .A2(_05451_),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11040_ (.A1(_05457_),
    .A2(_05450_),
    .B(_05458_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11041_ (.I(_01882_),
    .Z(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11042_ (.I(_05438_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11043_ (.I(_05440_),
    .Z(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11044_ (.A1(\as2650.stack[0][8] ),
    .A2(_05461_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11045_ (.A1(_05459_),
    .A2(_05460_),
    .B(_05462_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11046_ (.I(_01898_),
    .Z(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11047_ (.A1(\as2650.stack[0][9] ),
    .A2(_05461_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11048_ (.A1(_05463_),
    .A2(_05460_),
    .B(_05464_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11049_ (.I(_01912_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11050_ (.A1(\as2650.stack[0][10] ),
    .A2(_05461_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11051_ (.A1(_05465_),
    .A2(_05460_),
    .B(_05466_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11052_ (.I(_01927_),
    .Z(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11053_ (.A1(\as2650.stack[0][11] ),
    .A2(_05461_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11054_ (.A1(_05467_),
    .A2(_05460_),
    .B(_05468_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11055_ (.I(_01939_),
    .Z(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11056_ (.I(_05438_),
    .Z(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11057_ (.I(_05440_),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11058_ (.A1(\as2650.stack[0][12] ),
    .A2(_05471_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11059_ (.A1(_05469_),
    .A2(_05470_),
    .B(_05472_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11060_ (.I(_01946_),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11061_ (.A1(\as2650.stack[0][13] ),
    .A2(_05471_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11062_ (.A1(_05473_),
    .A2(_05470_),
    .B(_05474_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11063_ (.I(_01953_),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11064_ (.A1(\as2650.stack[0][14] ),
    .A2(_05471_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11065_ (.A1(_05475_),
    .A2(_05470_),
    .B(_05476_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11066_ (.I(_01958_),
    .Z(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11067_ (.A1(\as2650.stack[0][15] ),
    .A2(_05471_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11068_ (.A1(_05477_),
    .A2(_05470_),
    .B(_05478_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11069_ (.A1(_00180_),
    .A2(_01594_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11070_ (.A1(_04769_),
    .A2(_05142_),
    .A3(_04721_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11071_ (.I(_05479_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11072_ (.A1(_05168_),
    .A2(_05479_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11073_ (.I(_05481_),
    .Z(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11074_ (.I(\as2650.regs[7][0] ),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11075_ (.A1(_05163_),
    .A2(_05480_),
    .B1(_05482_),
    .B2(_05483_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11076_ (.I(\as2650.regs[7][1] ),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11077_ (.A1(_05171_),
    .A2(_05480_),
    .B1(_05482_),
    .B2(_05484_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11078_ (.I(\as2650.regs[7][2] ),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11079_ (.A1(_05172_),
    .A2(_05480_),
    .B1(_05482_),
    .B2(_05485_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11080_ (.I(\as2650.regs[7][3] ),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11081_ (.A1(_05173_),
    .A2(_05480_),
    .B1(_05482_),
    .B2(_05486_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11082_ (.I(_05479_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11083_ (.I(_05481_),
    .Z(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11084_ (.I(\as2650.regs[7][4] ),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11085_ (.A1(_05174_),
    .A2(_05487_),
    .B1(_05488_),
    .B2(_05489_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11086_ (.I(\as2650.regs[7][5] ),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11087_ (.A1(_05177_),
    .A2(_05487_),
    .B1(_05488_),
    .B2(_05490_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11088_ (.I(\as2650.regs[7][6] ),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11089_ (.A1(_05178_),
    .A2(_05487_),
    .B1(_05488_),
    .B2(_05491_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11090_ (.I(\as2650.regs[7][7] ),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11091_ (.A1(_05179_),
    .A2(_05487_),
    .B1(_05488_),
    .B2(_05492_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11092_ (.A1(_01685_),
    .A2(_05186_),
    .A3(_04622_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11093_ (.I(_05493_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11094_ (.I(_05494_),
    .Z(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11095_ (.I(_05493_),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11096_ (.I(_05496_),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11097_ (.A1(\as2650.stack[14][0] ),
    .A2(_05497_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11098_ (.A1(_05436_),
    .A2(_05495_),
    .B(_05498_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11099_ (.A1(\as2650.stack[14][1] ),
    .A2(_05497_),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11100_ (.A1(_05443_),
    .A2(_05495_),
    .B(_05499_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11101_ (.A1(\as2650.stack[14][2] ),
    .A2(_05497_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11102_ (.A1(_05445_),
    .A2(_05495_),
    .B(_05500_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11103_ (.A1(\as2650.stack[14][3] ),
    .A2(_05497_),
    .ZN(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11104_ (.A1(_05447_),
    .A2(_05495_),
    .B(_05501_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11105_ (.I(_05494_),
    .Z(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11106_ (.I(_05496_),
    .Z(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11107_ (.A1(\as2650.stack[14][4] ),
    .A2(_05503_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11108_ (.A1(_05449_),
    .A2(_05502_),
    .B(_05504_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11109_ (.A1(\as2650.stack[14][5] ),
    .A2(_05503_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11110_ (.A1(_05453_),
    .A2(_05502_),
    .B(_05505_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11111_ (.A1(\as2650.stack[14][6] ),
    .A2(_05503_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11112_ (.A1(_05455_),
    .A2(_05502_),
    .B(_05506_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11113_ (.A1(\as2650.stack[14][7] ),
    .A2(_05503_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11114_ (.A1(_05457_),
    .A2(_05502_),
    .B(_05507_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11115_ (.I(_05494_),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11116_ (.I(_05496_),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11117_ (.A1(\as2650.stack[14][8] ),
    .A2(_05509_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11118_ (.A1(_05459_),
    .A2(_05508_),
    .B(_05510_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11119_ (.A1(\as2650.stack[14][9] ),
    .A2(_05509_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11120_ (.A1(_05463_),
    .A2(_05508_),
    .B(_05511_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11121_ (.A1(\as2650.stack[14][10] ),
    .A2(_05509_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11122_ (.A1(_05465_),
    .A2(_05508_),
    .B(_05512_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11123_ (.A1(\as2650.stack[14][11] ),
    .A2(_05509_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11124_ (.A1(_05467_),
    .A2(_05508_),
    .B(_05513_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11125_ (.I(_05494_),
    .Z(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11126_ (.I(_05496_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11127_ (.A1(\as2650.stack[14][12] ),
    .A2(_05515_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11128_ (.A1(_05469_),
    .A2(_05514_),
    .B(_05516_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11129_ (.A1(\as2650.stack[14][13] ),
    .A2(_05515_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11130_ (.A1(_05473_),
    .A2(_05514_),
    .B(_05517_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11131_ (.A1(\as2650.stack[14][14] ),
    .A2(_05515_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11132_ (.A1(_05475_),
    .A2(_05514_),
    .B(_05518_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11133_ (.A1(\as2650.stack[14][15] ),
    .A2(_05515_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11134_ (.A1(_05477_),
    .A2(_05514_),
    .B(_05519_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11135_ (.A1(_01685_),
    .A2(_05186_),
    .A3(_04522_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11136_ (.I(_05520_),
    .Z(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11137_ (.I(_05521_),
    .Z(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11138_ (.I(_05520_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11139_ (.I(_05523_),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11140_ (.A1(\as2650.stack[13][0] ),
    .A2(_05524_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11141_ (.A1(_05436_),
    .A2(_05522_),
    .B(_05525_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11142_ (.A1(\as2650.stack[13][1] ),
    .A2(_05524_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11143_ (.A1(_05443_),
    .A2(_05522_),
    .B(_05526_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11144_ (.A1(\as2650.stack[13][2] ),
    .A2(_05524_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11145_ (.A1(_05445_),
    .A2(_05522_),
    .B(_05527_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11146_ (.A1(\as2650.stack[13][3] ),
    .A2(_05524_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11147_ (.A1(_05447_),
    .A2(_05522_),
    .B(_05528_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11148_ (.I(_05521_),
    .Z(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11149_ (.I(_05523_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11150_ (.A1(\as2650.stack[13][4] ),
    .A2(_05530_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11151_ (.A1(_05449_),
    .A2(_05529_),
    .B(_05531_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11152_ (.A1(\as2650.stack[13][5] ),
    .A2(_05530_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11153_ (.A1(_05453_),
    .A2(_05529_),
    .B(_05532_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11154_ (.A1(\as2650.stack[13][6] ),
    .A2(_05530_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11155_ (.A1(_05455_),
    .A2(_05529_),
    .B(_05533_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11156_ (.A1(\as2650.stack[13][7] ),
    .A2(_05530_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11157_ (.A1(_05457_),
    .A2(_05529_),
    .B(_05534_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11158_ (.I(_05521_),
    .Z(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11159_ (.I(_05523_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11160_ (.A1(\as2650.stack[13][8] ),
    .A2(_05536_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11161_ (.A1(_05459_),
    .A2(_05535_),
    .B(_05537_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11162_ (.A1(\as2650.stack[13][9] ),
    .A2(_05536_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11163_ (.A1(_05463_),
    .A2(_05535_),
    .B(_05538_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11164_ (.A1(\as2650.stack[13][10] ),
    .A2(_05536_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11165_ (.A1(_05465_),
    .A2(_05535_),
    .B(_05539_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11166_ (.A1(\as2650.stack[13][11] ),
    .A2(_05536_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11167_ (.A1(_05467_),
    .A2(_05535_),
    .B(_05540_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11168_ (.I(_05521_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11169_ (.I(_05523_),
    .Z(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11170_ (.A1(\as2650.stack[13][12] ),
    .A2(_05542_),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11171_ (.A1(_05469_),
    .A2(_05541_),
    .B(_05543_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11172_ (.A1(\as2650.stack[13][13] ),
    .A2(_05542_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11173_ (.A1(_05473_),
    .A2(_05541_),
    .B(_05544_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11174_ (.A1(\as2650.stack[13][14] ),
    .A2(_05542_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11175_ (.A1(_05475_),
    .A2(_05541_),
    .B(_05545_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11176_ (.A1(\as2650.stack[13][15] ),
    .A2(_05542_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11177_ (.A1(_05477_),
    .A2(_05541_),
    .B(_05546_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11178_ (.A1(_01713_),
    .A2(_01962_),
    .A3(_04522_),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11179_ (.I(_05547_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11180_ (.I(_05548_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11181_ (.I(_05547_),
    .Z(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11182_ (.I(_05550_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11183_ (.A1(\as2650.stack[9][0] ),
    .A2(_05551_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11184_ (.A1(_05436_),
    .A2(_05549_),
    .B(_05552_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11185_ (.A1(\as2650.stack[9][1] ),
    .A2(_05551_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11186_ (.A1(_05443_),
    .A2(_05549_),
    .B(_05553_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11187_ (.A1(\as2650.stack[9][2] ),
    .A2(_05551_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11188_ (.A1(_05445_),
    .A2(_05549_),
    .B(_05554_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11189_ (.A1(\as2650.stack[9][3] ),
    .A2(_05551_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11190_ (.A1(_05447_),
    .A2(_05549_),
    .B(_05555_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11191_ (.I(_05548_),
    .Z(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11192_ (.I(_05550_),
    .Z(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11193_ (.A1(\as2650.stack[9][4] ),
    .A2(_05557_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11194_ (.A1(_05449_),
    .A2(_05556_),
    .B(_05558_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11195_ (.A1(\as2650.stack[9][5] ),
    .A2(_05557_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11196_ (.A1(_05453_),
    .A2(_05556_),
    .B(_05559_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11197_ (.A1(\as2650.stack[9][6] ),
    .A2(_05557_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11198_ (.A1(_05455_),
    .A2(_05556_),
    .B(_05560_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11199_ (.A1(\as2650.stack[9][7] ),
    .A2(_05557_),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11200_ (.A1(_05457_),
    .A2(_05556_),
    .B(_05561_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11201_ (.I(_05548_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11202_ (.I(_05550_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11203_ (.A1(\as2650.stack[9][8] ),
    .A2(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11204_ (.A1(_05459_),
    .A2(_05562_),
    .B(_05564_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11205_ (.A1(\as2650.stack[9][9] ),
    .A2(_05563_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11206_ (.A1(_05463_),
    .A2(_05562_),
    .B(_05565_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11207_ (.A1(\as2650.stack[9][10] ),
    .A2(_05563_),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11208_ (.A1(_05465_),
    .A2(_05562_),
    .B(_05566_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11209_ (.A1(\as2650.stack[9][11] ),
    .A2(_05563_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11210_ (.A1(_05467_),
    .A2(_05562_),
    .B(_05567_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11211_ (.I(_05548_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11212_ (.I(_05550_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11213_ (.A1(\as2650.stack[9][12] ),
    .A2(_05569_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11214_ (.A1(_05469_),
    .A2(_05568_),
    .B(_05570_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11215_ (.A1(\as2650.stack[9][13] ),
    .A2(_05569_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11216_ (.A1(_05473_),
    .A2(_05568_),
    .B(_05571_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11217_ (.A1(\as2650.stack[9][14] ),
    .A2(_05569_),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11218_ (.A1(_05475_),
    .A2(_05568_),
    .B(_05572_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11219_ (.A1(\as2650.stack[9][15] ),
    .A2(_05569_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11220_ (.A1(_05477_),
    .A2(_05568_),
    .B(_05573_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11221_ (.D(_00017_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11222_ (.D(_00018_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11223_ (.D(_00019_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11224_ (.D(_00020_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11225_ (.D(_00021_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11226_ (.D(_00022_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11227_ (.D(_00023_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11228_ (.D(_00024_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11229_ (.D(_00025_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11230_ (.D(_00026_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11231_ (.D(_00027_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11232_ (.D(_00028_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11233_ (.D(_00029_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11234_ (.D(_00030_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11235_ (.D(_00031_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11236_ (.D(_00032_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11237_ (.D(_00033_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11238_ (.D(_00034_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11239_ (.D(_00035_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11240_ (.D(_00036_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11241_ (.D(_00037_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11242_ (.D(_00038_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11243_ (.D(_00039_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11244_ (.D(_00040_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11245_ (.D(_00041_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11246_ (.D(_00042_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11247_ (.D(_00043_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11248_ (.D(_00044_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11249_ (.D(_00045_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11250_ (.D(_00046_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11251_ (.D(_00047_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11252_ (.D(_00048_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11253_ (.D(_00049_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11254_ (.D(_00050_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(net122));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11255_ (.D(_00051_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(net129));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11256_ (.D(_00052_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(net130));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11257_ (.D(_00053_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(net131));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11258_ (.D(_00054_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11259_ (.D(_00055_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11260_ (.D(_00056_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11261_ (.D(_00057_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11262_ (.D(_00058_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11263_ (.D(_00059_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11264_ (.D(_00060_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(net123));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11265_ (.D(_00061_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(net124));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11266_ (.D(_00062_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(net125));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11267_ (.D(_00063_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(net126));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11268_ (.D(_00064_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net127));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11269_ (.D(_00065_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(net128));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11270_ (.D(_00066_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(net106));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11271_ (.D(_00067_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(net113));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11272_ (.D(_00068_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(net114));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11273_ (.D(_00069_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(net115));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11274_ (.D(_00070_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(net116));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11275_ (.D(_00071_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(net117));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11276_ (.D(_00072_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(net118));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11277_ (.D(_00073_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(net119));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11278_ (.D(_00074_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net120));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11279_ (.D(_00075_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net121));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11280_ (.D(_00076_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net107));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11281_ (.D(_00077_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(net108));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11282_ (.D(_00078_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(net109));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11283_ (.D(_00079_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(net110));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11284_ (.D(_00080_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(net111));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11285_ (.D(_00081_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(net112));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11286_ (.D(_00082_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(net239));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11287_ (.D(_00083_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(net159));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11288_ (.D(_00084_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(net160));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11289_ (.D(_00085_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(net161));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11290_ (.D(_00086_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net265));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11291_ (.D(_00087_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(net266));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11292_ (.D(_00088_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(net277));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11293_ (.D(_00089_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(net288));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11294_ (.D(_00090_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(net291));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11295_ (.D(_00091_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(net292));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11296_ (.D(_00092_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(net293));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11297_ (.D(_00093_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(net294));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11298_ (.D(_00094_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(net295));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11299_ (.D(_00095_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net296));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11300_ (.D(_00096_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net297));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11301_ (.D(_00097_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net267));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11302_ (.D(_00098_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(net268));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11303_ (.D(_00099_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(net269));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11304_ (.D(_00100_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(net270));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11305_ (.D(_00101_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(net271));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11306_ (.D(_00102_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(net272));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11307_ (.D(_00103_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(net273));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11308_ (.D(_00104_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net274));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11309_ (.D(_00105_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net275));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11310_ (.D(_00106_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(net276));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11311_ (.D(_00107_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net278));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11312_ (.D(_00108_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net279));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11313_ (.D(_00109_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net280));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11314_ (.D(_00110_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net281));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11315_ (.D(_00111_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(net282));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11316_ (.D(_00112_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net283));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11317_ (.D(_00113_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net284));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11318_ (.D(_00114_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(net285));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11319_ (.D(_00115_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(net286));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11320_ (.D(_00116_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(net287));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11321_ (.D(_00117_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(net289));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11322_ (.D(_00118_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(net290));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11323_ (.D(_00119_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11324_ (.D(_00120_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11325_ (.D(_00121_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(wb_debug_carry));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11326_ (.D(_00122_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\web_behavior[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11327_ (.D(net368),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\web_behavior[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11328_ (.D(net360),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(wb_reset_override_en));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11329_ (.D(net364),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(wb_reset_override));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11330_ (.D(net407),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(wb_io3_test));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11331_ (.D(net371),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(net182));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11332_ (.D(_00128_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11333_ (.D(_00129_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\wb_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11334_ (.D(_00130_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\wb_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11335_ (.D(_00131_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\wb_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11336_ (.D(_00132_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\wb_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11337_ (.D(_00133_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\wb_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11338_ (.D(_00134_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\wb_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11339_ (.D(_00135_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\wb_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11340_ (.D(_00136_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\wb_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11341_ (.D(_00137_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\wb_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11342_ (.D(_00138_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\wb_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11343_ (.D(net375),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\wb_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11344_ (.D(net379),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\wb_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11345_ (.D(_00141_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\wb_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11346_ (.D(_00142_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\wb_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11347_ (.D(_00143_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\wb_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11348_ (.D(_00144_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\wb_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11349_ (.D(_00145_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\wb_counter[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11350_ (.D(net383),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\wb_counter[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11351_ (.D(_00147_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\wb_counter[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11352_ (.D(_00148_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\wb_counter[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11353_ (.D(_00149_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\wb_counter[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11354_ (.D(_00150_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\wb_counter[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11355_ (.D(_00151_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\wb_counter[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11356_ (.D(_00152_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\wb_counter[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11357_ (.D(_00153_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\wb_counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11358_ (.D(_00154_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\wb_counter[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11359_ (.D(_00155_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\wb_counter[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11360_ (.D(_00156_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\wb_counter[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11361_ (.D(_00157_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\wb_counter[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11362_ (.D(_00158_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\wb_counter[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11363_ (.D(_00159_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\wb_counter[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11364_ (.D(_00160_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\wb_counter[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11365_ (.D(_00161_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net221));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11366_ (.D(_00162_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net228));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11367_ (.D(_00163_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net229));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11368_ (.D(_00164_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net230));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11369_ (.D(_00165_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net231));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11370_ (.D(_00166_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net232));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11371_ (.D(_00167_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net233));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11372_ (.D(_00168_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net234));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11373_ (.D(_00169_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11374_ (.D(_00170_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.insin[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11375_ (.D(_00171_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.insin[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11376_ (.D(_00172_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.insin[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11377_ (.D(_00173_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.insin[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11378_ (.D(_00174_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.insin[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11379_ (.D(_00175_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.insin[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11380_ (.D(_00176_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.indirect_target[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11381_ (.D(_00005_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11382_ (.D(_00008_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11383_ (.D(_00009_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11384_ (.D(_00010_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.is_interrupt_cycle ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11385_ (.D(_00011_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11386_ (.D(_00012_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11387_ (.D(_00013_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11388_ (.D(_00014_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11389_ (.D(_00015_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11390_ (.D(_00016_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11391_ (.D(_00006_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11392_ (.D(_00007_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11393_ (.D(_00177_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.cpu_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11394_ (.D(_00178_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.chirp_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11395_ (.D(_00179_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.chirp_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11396_ (.D(_00180_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.chirp_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11397_ (.D(_00181_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.indirect_target[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11398_ (.D(_00182_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.indirect_target[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11399_ (.D(_00183_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.indirect_target[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11400_ (.D(_00184_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.indirect_target[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11401_ (.D(_00185_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.indirect_target[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11402_ (.D(_00186_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.indirect_target[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11403_ (.D(_00187_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.indirect_target[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11404_ (.D(_00188_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.indirect_target[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11405_ (.D(_00189_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.indirect_target[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11406_ (.D(_00190_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.indirect_target[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11407_ (.D(_00191_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.indirect_target[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11408_ (.D(_00192_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.indirect_target[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11409_ (.D(_00193_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.indirect_target[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11410_ (.D(_00194_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.indirect_target[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11411_ (.D(_00195_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.indirect_target[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11412_ (.D(_00196_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.indexed_cyc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11413_ (.D(_00197_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.indexed_cyc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11414_ (.D(_00198_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.indirect_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11415_ (.D(_00199_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.extend ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11416_ (.D(_00200_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(net213));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11417_ (.D(_00201_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11418_ (.D(_00202_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11419_ (.D(_00203_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.instruction_args_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11420_ (.D(_00204_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11421_ (.D(_00205_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.instruction_args_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11422_ (.D(_00206_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11423_ (.D(_00207_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11424_ (.D(_00208_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.instruction_args_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11425_ (.D(_00209_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11426_ (.D(_00210_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11427_ (.D(_00211_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11428_ (.D(_00212_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11429_ (.D(_00213_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11430_ (.D(_00214_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11431_ (.D(_00215_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11432_ (.D(_00216_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.instruction_args_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11433_ (.D(_00217_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.instruction_args_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11434_ (.D(_00218_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11435_ (.D(_00219_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11436_ (.D(_00220_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11437_ (.D(_00221_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11438_ (.D(_00222_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11439_ (.D(_00223_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.insin[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11440_ (.D(_00224_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11441_ (.D(_00225_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11442_ (.D(_00226_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11443_ (.D(_00227_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11444_ (.D(_00228_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11445_ (.D(_00229_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11446_ (.D(_00230_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11447_ (.D(_00231_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11448_ (.D(_00232_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11449_ (.D(_00233_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.ivectors_base[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11450_ (.D(_00234_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.ivectors_base[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11451_ (.D(_00235_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11452_ (.D(_00236_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.PC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11453_ (.D(_00237_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11454_ (.D(_00238_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11455_ (.D(_00239_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.PC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11456_ (.D(_00240_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11457_ (.D(_00241_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11458_ (.D(_00242_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11459_ (.D(_00243_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11460_ (.D(_00244_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11461_ (.D(_00245_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11462_ (.D(_00246_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11463_ (.D(_00247_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11464_ (.D(_00248_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11465_ (.D(_00249_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.debug_psl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11466_ (.D(_00250_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11467_ (.D(_00251_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11468_ (.D(_00252_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11469_ (.D(_00253_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11470_ (.D(_00254_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.debug_psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11471_ (.D(_00255_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.debug_psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11472_ (.D(_00256_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11473_ (.D(_00257_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.debug_psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11474_ (.D(_00258_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.debug_psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11475_ (.D(_00259_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.debug_psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11476_ (.D(_00260_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11477_ (.D(_00261_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11478_ (.D(_00262_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(net181));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11479_ (.D(_00263_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11480_ (.D(_00264_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.irqs_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11481_ (.D(_00265_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.irqs_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11482_ (.D(_00266_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.irqs_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11483_ (.D(_00267_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.irqs_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11484_ (.D(_00268_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.irqs_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11485_ (.D(_00269_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.irqs_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11486_ (.D(_00270_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.irqs_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11487_ (.D(_00271_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11488_ (.D(_00272_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11489_ (.D(_00273_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11490_ (.D(_00274_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11491_ (.D(_00275_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11492_ (.D(_00276_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11493_ (.D(_00277_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11494_ (.D(_00278_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11495_ (.D(_00279_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11496_ (.D(_00280_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11497_ (.D(_00281_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11498_ (.D(_00282_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11499_ (.D(_00283_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11500_ (.D(_00284_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11501_ (.D(_00285_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11502_ (.D(_00286_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11503_ (.D(_00287_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11504_ (.D(_00288_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net147));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11505_ (.D(_00289_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net148));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11506_ (.D(_00290_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net149));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11507_ (.D(_00291_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net150));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11508_ (.D(_00292_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net151));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11509_ (.D(_00293_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net152));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11510_ (.D(_00294_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net153));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11511_ (.D(_00295_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net154));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11512_ (.D(_00296_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net146));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11513_ (.D(_00297_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(net140));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11514_ (.D(_00298_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(net141));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11515_ (.D(_00299_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(net142));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11516_ (.D(_00300_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(net143));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11517_ (.D(_00301_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11518_ (.D(_00302_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(net145));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11519_ (.D(_00303_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.ext_io_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11520_ (.D(_00304_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.ext_io_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11521_ (.D(_00305_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11522_ (.D(_00306_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net235));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11523_ (.D(_00307_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(net236));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11524_ (.D(_00308_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net222));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11525_ (.D(_00309_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net223));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11526_ (.D(_00310_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net224));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11527_ (.D(_00311_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net225));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11528_ (.D(_00312_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(net226));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11529_ (.D(_00313_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net227));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11530_ (.D(_00314_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11531_ (.D(_00315_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11532_ (.D(_00316_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11533_ (.D(_00317_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11534_ (.D(_00318_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11535_ (.D(_00319_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11536_ (.D(_00320_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11537_ (.D(_00321_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11538_ (.D(_00322_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11539_ (.D(_00323_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11540_ (.D(_00324_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11541_ (.D(_00325_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11542_ (.D(_00326_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11543_ (.D(_00327_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11544_ (.D(_00328_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11545_ (.D(_00329_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11546_ (.D(_00330_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11547_ (.D(_00331_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11548_ (.D(_00332_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11549_ (.D(_00333_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11550_ (.D(_00334_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11551_ (.D(_00335_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11552_ (.D(_00336_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11553_ (.D(_00337_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11554_ (.D(_00338_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11555_ (.D(_00339_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11556_ (.D(_00340_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11557_ (.D(_00341_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11558_ (.D(_00342_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11559_ (.D(_00343_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11560_ (.D(_00344_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11561_ (.D(_00345_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11562_ (.D(_00346_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11563_ (.D(_00347_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11564_ (.D(_00348_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11565_ (.D(_00349_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11566_ (.D(_00350_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11567_ (.D(_00351_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11568_ (.D(_00352_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11569_ (.D(_00353_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11570_ (.D(_00354_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11571_ (.D(_00355_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11572_ (.D(_00356_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11573_ (.D(_00357_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11574_ (.D(_00358_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11575_ (.D(_00359_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11576_ (.D(_00360_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11577_ (.D(_00361_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11578_ (.D(_00362_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11579_ (.D(_00363_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11580_ (.D(_00364_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11581_ (.D(_00365_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11582_ (.D(_00366_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11583_ (.D(_00367_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11584_ (.D(_00368_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11585_ (.D(_00369_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11586_ (.D(_00370_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11587_ (.D(_00371_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11588_ (.D(_00372_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11589_ (.D(_00373_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11590_ (.D(_00374_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11591_ (.D(_00375_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11592_ (.D(_00376_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11593_ (.D(_00377_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11594_ (.D(_00378_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11595_ (.D(_00379_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11596_ (.D(_00380_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11597_ (.D(_00381_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11598_ (.D(_00382_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11599_ (.D(_00383_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11600_ (.D(_00384_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11601_ (.D(_00385_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11602_ (.D(_00386_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11603_ (.D(_00387_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11604_ (.D(_00388_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11605_ (.D(_00389_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11606_ (.D(_00390_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11607_ (.D(_00391_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11608_ (.D(_00392_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11609_ (.D(_00393_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11610_ (.D(_00394_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11611_ (.D(_00395_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11612_ (.D(_00396_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11613_ (.D(_00397_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11614_ (.D(_00398_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11615_ (.D(_00399_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11616_ (.D(_00400_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11617_ (.D(_00401_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11618_ (.D(_00402_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11619_ (.D(_00403_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11620_ (.D(_00404_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11621_ (.D(_00405_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11622_ (.D(_00406_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11623_ (.D(_00407_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11624_ (.D(_00408_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11625_ (.D(_00409_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11626_ (.D(_00410_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11627_ (.D(_00411_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11628_ (.D(_00412_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11629_ (.D(_00413_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11630_ (.D(_00414_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11631_ (.D(_00415_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11632_ (.D(_00416_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11633_ (.D(_00417_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11634_ (.D(_00418_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11635_ (.D(_00419_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11636_ (.D(_00420_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11637_ (.D(_00421_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11638_ (.D(_00422_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11639_ (.D(_00423_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11640_ (.D(_00424_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11641_ (.D(_00425_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11642_ (.D(_00426_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11643_ (.D(_00427_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11644_ (.D(_00428_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11645_ (.D(_00429_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11646_ (.D(_00430_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11647_ (.D(_00431_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11648_ (.D(_00432_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11649_ (.D(_00433_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\as2650.stack[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11650_ (.D(_00434_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11651_ (.D(_00435_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11652_ (.D(_00436_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11653_ (.D(_00437_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11654_ (.D(_00438_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11655_ (.D(_00439_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11656_ (.D(_00440_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11657_ (.D(_00441_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11658_ (.D(_00442_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11659_ (.D(_00443_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11660_ (.D(_00444_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11661_ (.D(_00445_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11662_ (.D(_00446_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11663_ (.D(_00447_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11664_ (.D(_00448_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11665_ (.D(_00449_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11666_ (.D(_00450_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11667_ (.D(_00451_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11668_ (.D(_00452_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11669_ (.D(_00453_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11670_ (.D(_00454_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11671_ (.D(_00455_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11672_ (.D(_00456_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11673_ (.D(_00457_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.regs[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11674_ (.D(_00458_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11675_ (.D(_00459_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11676_ (.D(_00460_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11677_ (.D(_00461_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11678_ (.D(_00462_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11679_ (.D(_00463_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11680_ (.D(_00464_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11681_ (.D(_00465_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11682_ (.D(_00466_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11683_ (.D(_00467_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11684_ (.D(_00468_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00469_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00470_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00471_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00472_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00473_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00474_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.chirpchar[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00475_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00476_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00477_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00478_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00479_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00480_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11697_ (.D(_00481_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00482_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00483_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00484_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00485_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00486_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00487_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00488_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00489_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00490_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00491_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00492_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00493_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00494_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00495_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00496_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00497_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00498_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11715_ (.D(_00499_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00500_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00501_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00502_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00503_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00504_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00505_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00506_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00507_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11724_ (.D(_00508_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.regs[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00509_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00510_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00511_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00512_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00513_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00514_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00515_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00516_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00517_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00518_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00519_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00520_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00521_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00522_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00523_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00524_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00525_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00526_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00527_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00528_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00529_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00530_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00000_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.chirpchar[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00001_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.chirpchar[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00002_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.chirpchar[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00003_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.chirpchar[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00004_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.chirpchar[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00531_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.chirpchar[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00532_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00533_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00534_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00535_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00536_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00537_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00538_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00539_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11761_ (.D(_00540_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11762_ (.D(_00541_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11763_ (.D(_00542_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11764_ (.D(_00543_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11765_ (.D(_00544_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00545_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11767_ (.D(_00546_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11768_ (.D(_00547_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00548_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00549_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00550_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00551_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00552_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00553_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00554_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00555_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00556_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00557_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00558_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00559_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00560_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00561_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00562_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00563_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00564_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00565_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00566_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\as2650.stack[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00567_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00568_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00569_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00570_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00571_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00572_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00573_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00574_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00575_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00576_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00577_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00578_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00579_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00580_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00581_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00582_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00583_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00584_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00585_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00586_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00587_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11847_ (.I(net301),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11848_ (.I(net301),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11849_ (.I(net301),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11850_ (.I(net302),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11851_ (.I(net302),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11852_ (.I(net302),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11853_ (.I(net303),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11854_ (.I(net301),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11855_ (.I(net183),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11856_ (.I(net184),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11857_ (.I(net300),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11858_ (.I(net298),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11859_ (.I(net187),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11860_ (.I(net171),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11861_ (.I(net299),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11862_ (.I(net173),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0__01549_ (.I(_01549_),
    .Z(clknet_0__01549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f__01549_ (.I(clknet_0__01549_),
    .Z(clknet_1_0__leaf__01549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f__01549_ (.I(clknet_0__01549_),
    .Z(clknet_1_1__leaf__01549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_110_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_118_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_128_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_129_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_130_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_132_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_135_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_136_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_137_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_138_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_139_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_140_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_142_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_144_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_145_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_146_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_147_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_148_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_149_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_149_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_150_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_151_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_151_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_152_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_153_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_154_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_155_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_155_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_157_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout301 (.I(net302),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout302 (.I(net164),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout303 (.I(net164),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout306 (.I(net181),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold100 (.I(wbs_dat_i[21]),
    .Z(net446));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold101 (.I(wbs_dat_i[18]),
    .Z(net447));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold102 (.I(wbs_dat_i[14]),
    .Z(net448));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold103 (.I(wbs_dat_i[19]),
    .Z(net449));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold104 (.I(wbs_dat_i[8]),
    .Z(net450));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold105 (.I(wbs_dat_i[26]),
    .Z(net451));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold106 (.I(wbs_dat_i[15]),
    .Z(net452));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold107 (.I(wbs_dat_i[20]),
    .Z(net453));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold108 (.I(wbs_dat_i[25]),
    .Z(net454));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold109 (.I(wbs_dat_i[13]),
    .Z(net455));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold110 (.I(wbs_dat_i[30]),
    .Z(net456));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold111 (.I(wbs_dat_i[5]),
    .Z(net457));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold112 (.I(wbs_dat_i[24]),
    .Z(net458));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold113 (.I(wbs_dat_i[2]),
    .Z(net459));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold114 (.I(wbs_adr_i[21]),
    .Z(net460));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold115 (.I(wbs_dat_i[0]),
    .Z(net461));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold116 (.I(wbs_dat_i[17]),
    .Z(net462));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold117 (.I(wbs_dat_i[16]),
    .Z(net463));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold118 (.I(wbs_dat_i[1]),
    .Z(net464));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold119 (.I(wbs_dat_i[23]),
    .Z(net465));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold120 (.I(wbs_stb_i),
    .Z(net466));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold121 (.I(wbs_dat_i[22]),
    .Z(net467));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(net435),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(net98),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(_02311_),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(_00124_),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(net457),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold18 (.I(net99),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(_02313_),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(_00125_),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(net432),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold22 (.I(net97),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(_02308_),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(_00123_),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(net431),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(_02316_),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(_00127_),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(wbs_dat_i[10]),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(net73),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(_02366_),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(_00139_),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(net440),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(net74),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(_02369_),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(_00140_),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(net462),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(net80),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(_02395_),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(_00146_),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(net444),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(net463),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(net79),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(net441),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(net75),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(net445),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(net100),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(net438),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold48 (.I(net93),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(net450),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(net102),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(net455),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(net76),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(net448),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(net77),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(net456),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold56 (.I(net95),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(net452),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(net78),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(net442),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(net103),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(net434),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(net460),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(_00126_),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(net436),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(_02028_),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(wbs_adr_i[20]),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(_02068_),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(net447),
    .Z(net412));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(net449),
    .Z(net413));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(net453),
    .Z(net414));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(net439),
    .Z(net415));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(net459),
    .Z(net416));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(net443),
    .Z(net417));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(net464),
    .Z(net418));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(net446),
    .Z(net419));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(net461),
    .Z(net420));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(net454),
    .Z(net421));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(net451),
    .Z(net422));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(net465),
    .Z(net423));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(net458),
    .Z(net424));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(net467),
    .Z(net425));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(wbs_cyc_i),
    .Z(net426));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold83 (.I(_02005_),
    .Z(net427));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(wbs_we_i),
    .Z(net428));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold85 (.I(wbs_dat_i[7]),
    .Z(net431));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold86 (.I(wbs_dat_i[3]),
    .Z(net432));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold87 (.I(_02334_),
    .Z(net433));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold88 (.I(wbs_dat_i[31]),
    .Z(net434));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold89 (.I(wbs_dat_i[4]),
    .Z(net435));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold90 (.I(wbs_adr_i[19]),
    .Z(net436));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold91 (.I(_02068_),
    .Z(net437));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold92 (.I(wbs_dat_i[29]),
    .Z(net438));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold93 (.I(wbs_dat_i[27]),
    .Z(net439));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold94 (.I(wbs_dat_i[11]),
    .Z(net440));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold95 (.I(wbs_dat_i[12]),
    .Z(net441));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold96 (.I(wbs_dat_i[9]),
    .Z(net442));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold97 (.I(wbs_dat_i[28]),
    .Z(net443));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold98 (.I(wbs_adr_i[22]),
    .Z(net444));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold99 (.I(wbs_dat_i[6]),
    .Z(net445));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(bus_in_gpios[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(bus_in_serial_ports[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input100 (.I(net389),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input101 (.I(net369),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input102 (.I(net393),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input103 (.I(net403),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input104 (.I(net466),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input105 (.I(net428),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(bus_in_serial_ports[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(bus_in_serial_ports[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(bus_in_serial_ports[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input14 (.I(bus_in_serial_ports[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(bus_in_serial_ports[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(bus_in_serial_ports[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(bus_in_sid[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(bus_in_sid[1]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(bus_in_sid[2]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(bus_in_gpios[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(bus_in_sid[3]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(bus_in_sid[4]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(bus_in_sid[5]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(bus_in_sid[6]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(bus_in_sid[7]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(bus_in_timers[0]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(bus_in_timers[1]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(bus_in_timers[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(bus_in_timers[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(bus_in_timers[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(bus_in_gpios[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(bus_in_timers[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(bus_in_timers[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(bus_in_timers[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input33 (.I(io_in[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(io_in[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(io_in[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(io_in[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input37 (.I(io_in[4]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(io_in[5]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(io_in[6]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(bus_in_gpios[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(io_in[7]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(io_in[8]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(io_in[9]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input43 (.I(irqs[0]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input44 (.I(irqs[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input45 (.I(irqs[2]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(irqs[3]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(irqs[4]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(irqs[5]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(irqs[6]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(bus_in_gpios[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(ram_bus_in[0]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(ram_bus_in[1]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(ram_bus_in[2]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(ram_bus_in[3]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(ram_bus_in[4]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(ram_bus_in[5]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(ram_bus_in[6]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(ram_bus_in[7]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input58 (.I(rom_bus_in[0]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input59 (.I(rom_bus_in[1]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(bus_in_gpios[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input60 (.I(rom_bus_in[2]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input61 (.I(rom_bus_in[3]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input62 (.I(rom_bus_in[4]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input63 (.I(rom_bus_in[5]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input64 (.I(rom_bus_in[6]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input65 (.I(rom_bus_in[7]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input66 (.I(wb_rst_i),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input67 (.I(net408),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input68 (.I(net410),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input69 (.I(net406),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(bus_in_gpios[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input70 (.I(net384),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(net426),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input72 (.I(net420),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input73 (.I(net372),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input74 (.I(net376),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input75 (.I(net387),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(net395),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(net397),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(net401),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(net385),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(bus_in_gpios[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(net380),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input81 (.I(net412),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input82 (.I(net413),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input83 (.I(net418),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input84 (.I(net414),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input85 (.I(net419),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input86 (.I(net425),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input87 (.I(net423),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input88 (.I(net424),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input89 (.I(net421),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(bus_in_serial_ports[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input90 (.I(net422),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input91 (.I(net415),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input92 (.I(net417),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input93 (.I(net391),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input94 (.I(net416),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input95 (.I(net399),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input96 (.I(net405),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input97 (.I(net365),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input98 (.I(net357),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input99 (.I(net361),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap304 (.I(_01535_),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap305 (.I(_00608_),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(RAM_end_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(RAM_end_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(RAM_end_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(RAM_end_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(RAM_end_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(RAM_end_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(RAM_end_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(RAM_end_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(RAM_end_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(RAM_end_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(RAM_end_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(RAM_end_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(RAM_end_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(RAM_end_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(RAM_end_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(RAM_end_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(RAM_start_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(RAM_start_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output124 (.I(net124),
    .Z(RAM_start_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output125 (.I(net125),
    .Z(RAM_start_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output126 (.I(net126),
    .Z(RAM_start_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output127 (.I(net127),
    .Z(RAM_start_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output128 (.I(net128),
    .Z(RAM_start_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output129 (.I(net129),
    .Z(RAM_start_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output130 (.I(net130),
    .Z(RAM_start_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output131 (.I(net131),
    .Z(RAM_start_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output132 (.I(net132),
    .Z(RAM_start_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output133 (.I(net133),
    .Z(RAM_start_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output134 (.I(net134),
    .Z(RAM_start_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output135 (.I(net135),
    .Z(RAM_start_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output136 (.I(net136),
    .Z(RAM_start_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output137 (.I(net137),
    .Z(RAM_start_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output138 (.I(net138),
    .Z(WEb_ram));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output139 (.I(net139),
    .Z(boot_rom_en));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output140 (.I(net140),
    .Z(bus_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output141 (.I(net141),
    .Z(bus_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output142 (.I(net142),
    .Z(bus_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output143 (.I(net143),
    .Z(bus_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output144 (.I(net144),
    .Z(bus_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output145 (.I(net145),
    .Z(bus_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output146 (.I(net146),
    .Z(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output147 (.I(net147),
    .Z(bus_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output148 (.I(net148),
    .Z(bus_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output149 (.I(net149),
    .Z(bus_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output150 (.I(net150),
    .Z(bus_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output151 (.I(net151),
    .Z(bus_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output152 (.I(net152),
    .Z(bus_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output153 (.I(net153),
    .Z(bus_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output154 (.I(net154),
    .Z(bus_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output155 (.I(net155),
    .Z(bus_we_gpios));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output156 (.I(net156),
    .Z(bus_we_serial_ports));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output157 (.I(net157),
    .Z(bus_we_sid));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output158 (.I(net158),
    .Z(bus_we_timers));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output159 (.I(net159),
    .Z(cs_port[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output160 (.I(net160),
    .Z(cs_port[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output161 (.I(net161),
    .Z(cs_port[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output162 (.I(net162),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output163 (.I(net163),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output164 (.I(net303),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output165 (.I(net165),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output166 (.I(net166),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output167 (.I(net167),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output168 (.I(net168),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output169 (.I(net169),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output170 (.I(net170),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output171 (.I(net171),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output172 (.I(net299),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output173 (.I(net173),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output174 (.I(net174),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output175 (.I(net175),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output176 (.I(net176),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output177 (.I(net177),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output178 (.I(net178),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output179 (.I(net179),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output180 (.I(net180),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output181 (.I(net306),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output182 (.I(net182),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output183 (.I(net183),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output184 (.I(net184),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output185 (.I(net300),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output186 (.I(net298),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output187 (.I(net187),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output188 (.I(net188),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output189 (.I(net189),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output190 (.I(net190),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output191 (.I(net191),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output192 (.I(net192),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output193 (.I(net193),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output194 (.I(net194),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output195 (.I(net195),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output196 (.I(net196),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output197 (.I(net197),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output198 (.I(net198),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output199 (.I(net199),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output200 (.I(net200),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output201 (.I(net201),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output202 (.I(net202),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output203 (.I(net203),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output204 (.I(net204),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output205 (.I(net205),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output206 (.I(net206),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output207 (.I(net207),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output208 (.I(net208),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output209 (.I(net209),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output210 (.I(net210),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output211 (.I(net211),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output212 (.I(net212),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output213 (.I(net213),
    .Z(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output214 (.I(net214),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output215 (.I(net215),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output216 (.I(net216),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output217 (.I(net217),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output218 (.I(net218),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output219 (.I(net219),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output220 (.I(net220),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output221 (.I(net221),
    .Z(last_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output222 (.I(net222),
    .Z(last_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output223 (.I(net223),
    .Z(last_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output224 (.I(net224),
    .Z(last_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output225 (.I(net225),
    .Z(last_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output226 (.I(net226),
    .Z(last_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output227 (.I(net227),
    .Z(last_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output228 (.I(net228),
    .Z(last_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output229 (.I(net229),
    .Z(last_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output230 (.I(net230),
    .Z(last_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output231 (.I(net231),
    .Z(last_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output232 (.I(net232),
    .Z(last_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output233 (.I(net233),
    .Z(last_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output234 (.I(net234),
    .Z(last_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output235 (.I(net235),
    .Z(last_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output236 (.I(net236),
    .Z(last_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output237 (.I(net237),
    .Z(le_hi_act));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output238 (.I(net238),
    .Z(le_lo_act));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output239 (.I(net239),
    .Z(ram_enabled));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output240 (.I(net240),
    .Z(requested_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output241 (.I(net241),
    .Z(requested_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output242 (.I(net242),
    .Z(requested_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output243 (.I(net243),
    .Z(requested_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output244 (.I(net244),
    .Z(requested_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output245 (.I(net245),
    .Z(requested_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output246 (.I(net246),
    .Z(requested_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output247 (.I(net247),
    .Z(requested_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output248 (.I(net248),
    .Z(requested_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output249 (.I(net249),
    .Z(requested_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output250 (.I(net250),
    .Z(requested_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output251 (.I(net251),
    .Z(requested_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output252 (.I(net252),
    .Z(requested_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output253 (.I(net253),
    .Z(requested_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output254 (.I(net254),
    .Z(requested_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output255 (.I(net255),
    .Z(requested_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output256 (.I(net355),
    .Z(reset_out));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output257 (.I(net257),
    .Z(rom_bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output258 (.I(net258),
    .Z(rom_bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output259 (.I(net259),
    .Z(rom_bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output260 (.I(net260),
    .Z(rom_bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output261 (.I(net261),
    .Z(rom_bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output262 (.I(net262),
    .Z(rom_bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output263 (.I(net263),
    .Z(rom_bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output264 (.I(net264),
    .Z(rom_bus_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output265 (.I(net265),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output266 (.I(net266),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output267 (.I(net267),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output268 (.I(net268),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output269 (.I(net269),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output270 (.I(net270),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output271 (.I(net271),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output272 (.I(net272),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output273 (.I(net273),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output274 (.I(net274),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output275 (.I(net275),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output276 (.I(net276),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output277 (.I(net277),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output278 (.I(net278),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output279 (.I(net279),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output280 (.I(net280),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output281 (.I(net281),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output282 (.I(net282),
    .Z(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output283 (.I(net283),
    .Z(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output284 (.I(net284),
    .Z(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output285 (.I(net285),
    .Z(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output286 (.I(net286),
    .Z(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output287 (.I(net287),
    .Z(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output288 (.I(net288),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output289 (.I(net289),
    .Z(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output290 (.I(net290),
    .Z(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output291 (.I(net291),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output292 (.I(net292),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output293 (.I(net293),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output294 (.I(net294),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output295 (.I(net295),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output296 (.I(net296),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output297 (.I(net297),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 rebuffer1 (.I(_00733_),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer10 (.I(_04059_),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 rebuffer11 (.I(net256),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(_01357_),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer13 (.I(_00938_),
    .Z(net429));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer14 (.I(_00619_),
    .Z(net430));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer2 (.I(net345),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer3 (.I(_00924_),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer4 (.I(_00934_),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(net352),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer6 (.I(net349),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer7 (.I(_01072_),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer8 (.I(_00907_),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 rebuffer9 (.I(_00906_),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire298 (.I(net186),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire299 (.I(net172),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire300 (.I(net185),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_307 (.ZN(net307));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_308 (.ZN(net308));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_309 (.ZN(net309));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_310 (.ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_311 (.ZN(net311));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_312 (.ZN(net312));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_313 (.ZN(net313));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_314 (.ZN(net314));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_315 (.ZN(net315));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_316 (.ZN(net316));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_317 (.ZN(net317));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_318 (.ZN(net318));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_319 (.ZN(net319));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_320 (.ZN(net320));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_321 (.ZN(net321));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_322 (.ZN(net322));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_323 (.ZN(net323));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_324 (.ZN(net324));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_325 (.ZN(net325));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_326 (.ZN(net326));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_327 (.ZN(net327));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_328 (.Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_329 (.Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_330 (.Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_331 (.Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_332 (.Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_333 (.Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_334 (.Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_335 (.Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_336 (.Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_337 (.Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_338 (.Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_339 (.Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_340 (.Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_341 (.Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_342 (.Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_343 (.Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_344 (.Z(net344));
 assign io_oeb[0] = net328;
 assign io_oeb[13] = net309;
 assign io_oeb[14] = net310;
 assign io_oeb[15] = net311;
 assign io_oeb[16] = net312;
 assign io_oeb[17] = net313;
 assign io_oeb[18] = net314;
 assign io_oeb[1] = net307;
 assign io_oeb[2] = net308;
 assign io_oeb[4] = net329;
 assign io_out[0] = net315;
 assign io_out[4] = net316;
 assign irq[0] = net317;
 assign irq[1] = net318;
 assign irq[2] = net319;
 assign la_data_out[33] = net330;
 assign la_data_out[34] = net331;
 assign la_data_out[35] = net332;
 assign la_data_out[36] = net333;
 assign la_data_out[37] = net334;
 assign la_data_out[38] = net335;
 assign la_data_out[39] = net336;
 assign la_data_out[40] = net337;
 assign la_data_out[41] = net320;
 assign la_data_out[42] = net321;
 assign la_data_out[43] = net322;
 assign la_data_out[44] = net323;
 assign la_data_out[45] = net324;
 assign la_data_out[46] = net325;
 assign la_data_out[47] = net326;
 assign la_data_out[48] = net327;
 assign la_data_out[49] = net338;
 assign la_data_out[50] = net339;
 assign la_data_out[51] = net340;
 assign la_data_out[52] = net341;
 assign la_data_out[53] = net342;
 assign la_data_out[54] = net343;
 assign la_data_out[55] = net344;
endmodule

