VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as2650
  CLASS BLOCK ;
  FOREIGN wrapped_as2650 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 750.000 ;
  PIN RAM_end_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 434.560 4.000 435.120 ;
    END
  END RAM_end_addr[0]
  PIN RAM_end_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 501.760 4.000 502.320 ;
    END
  END RAM_end_addr[10]
  PIN RAM_end_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 508.480 4.000 509.040 ;
    END
  END RAM_end_addr[11]
  PIN RAM_end_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 515.200 4.000 515.760 ;
    END
  END RAM_end_addr[12]
  PIN RAM_end_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.920 4.000 522.480 ;
    END
  END RAM_end_addr[13]
  PIN RAM_end_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 528.640 4.000 529.200 ;
    END
  END RAM_end_addr[14]
  PIN RAM_end_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 535.360 4.000 535.920 ;
    END
  END RAM_end_addr[15]
  PIN RAM_end_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 441.280 4.000 441.840 ;
    END
  END RAM_end_addr[1]
  PIN RAM_end_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END RAM_end_addr[2]
  PIN RAM_end_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.720 4.000 455.280 ;
    END
  END RAM_end_addr[3]
  PIN RAM_end_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 461.440 4.000 462.000 ;
    END
  END RAM_end_addr[4]
  PIN RAM_end_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 468.160 4.000 468.720 ;
    END
  END RAM_end_addr[5]
  PIN RAM_end_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 474.880 4.000 475.440 ;
    END
  END RAM_end_addr[6]
  PIN RAM_end_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 481.600 4.000 482.160 ;
    END
  END RAM_end_addr[7]
  PIN RAM_end_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 488.320 4.000 488.880 ;
    END
  END RAM_end_addr[8]
  PIN RAM_end_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 495.040 4.000 495.600 ;
    END
  END RAM_end_addr[9]
  PIN RAM_start_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 300.160 4.000 300.720 ;
    END
  END RAM_start_addr[0]
  PIN RAM_start_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 367.360 4.000 367.920 ;
    END
  END RAM_start_addr[10]
  PIN RAM_start_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.080 4.000 374.640 ;
    END
  END RAM_start_addr[11]
  PIN RAM_start_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END RAM_start_addr[12]
  PIN RAM_start_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 387.520 4.000 388.080 ;
    END
  END RAM_start_addr[13]
  PIN RAM_start_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 394.240 4.000 394.800 ;
    END
  END RAM_start_addr[14]
  PIN RAM_start_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 400.960 4.000 401.520 ;
    END
  END RAM_start_addr[15]
  PIN RAM_start_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.880 4.000 307.440 ;
    END
  END RAM_start_addr[1]
  PIN RAM_start_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.600 4.000 314.160 ;
    END
  END RAM_start_addr[2]
  PIN RAM_start_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 320.320 4.000 320.880 ;
    END
  END RAM_start_addr[3]
  PIN RAM_start_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 327.040 4.000 327.600 ;
    END
  END RAM_start_addr[4]
  PIN RAM_start_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 333.760 4.000 334.320 ;
    END
  END RAM_start_addr[5]
  PIN RAM_start_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 340.480 4.000 341.040 ;
    END
  END RAM_start_addr[6]
  PIN RAM_start_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.200 4.000 347.760 ;
    END
  END RAM_start_addr[7]
  PIN RAM_start_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 353.920 4.000 354.480 ;
    END
  END RAM_start_addr[8]
  PIN RAM_start_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 360.640 4.000 361.200 ;
    END
  END RAM_start_addr[9]
  PIN WEb_raw
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1022.560 746.000 1023.120 750.000 ;
    END
  END WEb_raw
  PIN boot_rom_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 427.840 4.000 428.400 ;
    END
  END boot_rom_en
  PIN bus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 746.000 740.880 750.000 ;
    END
  END bus_addr[0]
  PIN bus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 746.000 761.040 750.000 ;
    END
  END bus_addr[1]
  PIN bus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 780.640 746.000 781.200 750.000 ;
    END
  END bus_addr[2]
  PIN bus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 800.800 746.000 801.360 750.000 ;
    END
  END bus_addr[3]
  PIN bus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 820.960 746.000 821.520 750.000 ;
    END
  END bus_addr[4]
  PIN bus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 841.120 746.000 841.680 750.000 ;
    END
  END bus_addr[5]
  PIN bus_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 720.160 746.000 720.720 750.000 ;
    END
  END bus_cyc
  PIN bus_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 746.000 559.440 750.000 ;
    END
  END bus_data_out[0]
  PIN bus_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 746.000 579.600 750.000 ;
    END
  END bus_data_out[1]
  PIN bus_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 746.000 599.760 750.000 ;
    END
  END bus_data_out[2]
  PIN bus_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 619.360 746.000 619.920 750.000 ;
    END
  END bus_data_out[3]
  PIN bus_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 746.000 640.080 750.000 ;
    END
  END bus_data_out[4]
  PIN bus_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 746.000 660.240 750.000 ;
    END
  END bus_data_out[5]
  PIN bus_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 679.840 746.000 680.400 750.000 ;
    END
  END bus_data_out[6]
  PIN bus_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 700.000 746.000 700.560 750.000 ;
    END
  END bus_data_out[7]
  PIN bus_in_gpios[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 431.200 1100.000 431.760 ;
    END
  END bus_in_gpios[0]
  PIN bus_in_gpios[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 437.920 1100.000 438.480 ;
    END
  END bus_in_gpios[1]
  PIN bus_in_gpios[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 444.640 1100.000 445.200 ;
    END
  END bus_in_gpios[2]
  PIN bus_in_gpios[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 451.360 1100.000 451.920 ;
    END
  END bus_in_gpios[3]
  PIN bus_in_gpios[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 458.080 1100.000 458.640 ;
    END
  END bus_in_gpios[4]
  PIN bus_in_gpios[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 464.800 1100.000 465.360 ;
    END
  END bus_in_gpios[5]
  PIN bus_in_gpios[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 471.520 1100.000 472.080 ;
    END
  END bus_in_gpios[6]
  PIN bus_in_gpios[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 478.240 1100.000 478.800 ;
    END
  END bus_in_gpios[7]
  PIN bus_in_serial_ports[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 746.000 861.840 750.000 ;
    END
  END bus_in_serial_ports[0]
  PIN bus_in_serial_ports[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 881.440 746.000 882.000 750.000 ;
    END
  END bus_in_serial_ports[1]
  PIN bus_in_serial_ports[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 901.600 746.000 902.160 750.000 ;
    END
  END bus_in_serial_ports[2]
  PIN bus_in_serial_ports[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 921.760 746.000 922.320 750.000 ;
    END
  END bus_in_serial_ports[3]
  PIN bus_in_serial_ports[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 941.920 746.000 942.480 750.000 ;
    END
  END bus_in_serial_ports[4]
  PIN bus_in_serial_ports[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 962.080 746.000 962.640 750.000 ;
    END
  END bus_in_serial_ports[5]
  PIN bus_in_serial_ports[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 982.240 746.000 982.800 750.000 ;
    END
  END bus_in_serial_ports[6]
  PIN bus_in_serial_ports[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1002.400 746.000 1002.960 750.000 ;
    END
  END bus_in_serial_ports[7]
  PIN bus_in_sid[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 565.600 1100.000 566.160 ;
    END
  END bus_in_sid[0]
  PIN bus_in_sid[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 572.320 1100.000 572.880 ;
    END
  END bus_in_sid[1]
  PIN bus_in_sid[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 579.040 1100.000 579.600 ;
    END
  END bus_in_sid[2]
  PIN bus_in_sid[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 585.760 1100.000 586.320 ;
    END
  END bus_in_sid[3]
  PIN bus_in_sid[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 592.480 1100.000 593.040 ;
    END
  END bus_in_sid[4]
  PIN bus_in_sid[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 599.200 1100.000 599.760 ;
    END
  END bus_in_sid[5]
  PIN bus_in_sid[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 605.920 1100.000 606.480 ;
    END
  END bus_in_sid[6]
  PIN bus_in_sid[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 612.640 1100.000 613.200 ;
    END
  END bus_in_sid[7]
  PIN bus_in_timers[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 505.120 1100.000 505.680 ;
    END
  END bus_in_timers[0]
  PIN bus_in_timers[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 511.840 1100.000 512.400 ;
    END
  END bus_in_timers[1]
  PIN bus_in_timers[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 518.560 1100.000 519.120 ;
    END
  END bus_in_timers[2]
  PIN bus_in_timers[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 525.280 1100.000 525.840 ;
    END
  END bus_in_timers[3]
  PIN bus_in_timers[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 532.000 1100.000 532.560 ;
    END
  END bus_in_timers[4]
  PIN bus_in_timers[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 538.720 1100.000 539.280 ;
    END
  END bus_in_timers[5]
  PIN bus_in_timers[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 545.440 1100.000 546.000 ;
    END
  END bus_in_timers[6]
  PIN bus_in_timers[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 552.160 1100.000 552.720 ;
    END
  END bus_in_timers[7]
  PIN bus_we_gpios
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 424.480 1100.000 425.040 ;
    END
  END bus_we_gpios
  PIN bus_we_serial_ports
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 498.400 1100.000 498.960 ;
    END
  END bus_we_serial_ports
  PIN bus_we_sid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 558.880 1100.000 559.440 ;
    END
  END bus_we_sid
  PIN bus_we_timers
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 491.680 1100.000 492.240 ;
    END
  END bus_we_timers
  PIN cs_port[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 407.680 4.000 408.240 ;
    END
  END cs_port[0]
  PIN cs_port[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 414.400 4.000 414.960 ;
    END
  END cs_port[1]
  PIN cs_port[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 421.120 4.000 421.680 ;
    END
  END cs_port[2]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 746.000 35.280 750.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 746.000 236.880 750.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 746.000 257.040 750.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 746.000 277.200 750.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 746.000 297.360 750.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 746.000 317.520 750.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 746.000 337.680 750.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 746.000 357.840 750.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 746.000 378.000 750.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 746.000 398.160 750.000 ;
    END
  END io_in[18]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 746.000 55.440 750.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 746.000 75.600 750.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 746.000 95.760 750.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 746.000 115.920 750.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 746.000 136.080 750.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 746.000 156.240 750.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 746.000 176.400 750.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 746.000 196.560 750.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 746.000 216.720 750.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 172.480 4.000 173.040 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 239.680 4.000 240.240 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.400 4.000 246.960 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.120 4.000 253.680 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 259.840 4.000 260.400 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.560 4.000 267.120 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 273.280 4.000 273.840 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.000 4.000 280.560 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.720 4.000 287.280 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 293.440 4.000 294.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.200 4.000 179.760 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 4.000 186.480 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 192.640 4.000 193.200 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 4.000 199.920 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.080 4.000 206.640 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 219.520 4.000 220.080 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.240 4.000 226.800 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.960 4.000 233.520 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.800 4.000 45.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.000 4.000 112.560 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 125.440 4.000 126.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 4.000 132.720 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 138.880 4.000 139.440 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.600 4.000 146.160 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.040 4.000 159.600 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 165.760 4.000 166.320 ;
    END
  END io_out[18]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 4.000 52.080 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.240 4.000 58.800 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.960 4.000 65.520 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 71.680 4.000 72.240 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.120 4.000 85.680 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 91.840 4.000 92.400 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 98.560 4.000 99.120 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 404.320 1100.000 404.880 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 411.040 1100.000 411.600 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 417.760 1100.000 418.320 ;
    END
  END irq[2]
  PIN irqs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 746.000 418.320 750.000 ;
    END
  END irqs[0]
  PIN irqs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 746.000 438.480 750.000 ;
    END
  END irqs[1]
  PIN irqs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 746.000 458.640 750.000 ;
    END
  END irqs[2]
  PIN irqs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 746.000 478.800 750.000 ;
    END
  END irqs[3]
  PIN irqs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 746.000 498.960 750.000 ;
    END
  END irqs[4]
  PIN irqs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 518.560 746.000 519.120 750.000 ;
    END
  END irqs[5]
  PIN irqs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 746.000 539.280 750.000 ;
    END
  END irqs[6]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 28.000 1100.000 28.560 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 95.200 1100.000 95.760 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 101.920 1100.000 102.480 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 108.640 1100.000 109.200 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 115.360 1100.000 115.920 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 122.080 1100.000 122.640 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 128.800 1100.000 129.360 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 135.520 1100.000 136.080 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 142.240 1100.000 142.800 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 148.960 1100.000 149.520 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 155.680 1100.000 156.240 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 34.720 1100.000 35.280 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 162.400 1100.000 162.960 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 169.120 1100.000 169.680 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 175.840 1100.000 176.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 182.560 1100.000 183.120 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 189.280 1100.000 189.840 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 196.000 1100.000 196.560 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 202.720 1100.000 203.280 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 209.440 1100.000 210.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 216.160 1100.000 216.720 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 222.880 1100.000 223.440 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 41.440 1100.000 42.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 229.600 1100.000 230.160 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 236.320 1100.000 236.880 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 243.040 1100.000 243.600 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 249.760 1100.000 250.320 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 256.480 1100.000 257.040 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 263.200 1100.000 263.760 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 269.920 1100.000 270.480 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 276.640 1100.000 277.200 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 283.360 1100.000 283.920 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 290.080 1100.000 290.640 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 48.160 1100.000 48.720 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 296.800 1100.000 297.360 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 303.520 1100.000 304.080 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 310.240 1100.000 310.800 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 316.960 1100.000 317.520 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 323.680 1100.000 324.240 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 330.400 1100.000 330.960 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 337.120 1100.000 337.680 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 343.840 1100.000 344.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 350.560 1100.000 351.120 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 357.280 1100.000 357.840 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 54.880 1100.000 55.440 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 364.000 1100.000 364.560 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 370.720 1100.000 371.280 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 377.440 1100.000 378.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 384.160 1100.000 384.720 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 390.880 1100.000 391.440 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 397.600 1100.000 398.160 ;
    END
  END la_data_out[55]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 61.600 1100.000 62.160 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 68.320 1100.000 68.880 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 75.040 1100.000 75.600 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 81.760 1100.000 82.320 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 88.480 1100.000 89.040 ;
    END
  END la_data_out[9]
  PIN last_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 938.560 0.000 939.120 4.000 ;
    END
  END last_addr[0]
  PIN last_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 0.000 1028.720 4.000 ;
    END
  END last_addr[10]
  PIN last_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1037.120 0.000 1037.680 4.000 ;
    END
  END last_addr[11]
  PIN last_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1046.080 0.000 1046.640 4.000 ;
    END
  END last_addr[12]
  PIN last_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 0.000 1055.600 4.000 ;
    END
  END last_addr[13]
  PIN last_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1064.000 0.000 1064.560 4.000 ;
    END
  END last_addr[14]
  PIN last_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1072.960 0.000 1073.520 4.000 ;
    END
  END last_addr[15]
  PIN last_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 0.000 948.080 4.000 ;
    END
  END last_addr[1]
  PIN last_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 956.480 0.000 957.040 4.000 ;
    END
  END last_addr[2]
  PIN last_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 965.440 0.000 966.000 4.000 ;
    END
  END last_addr[3]
  PIN last_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 0.000 974.960 4.000 ;
    END
  END last_addr[4]
  PIN last_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 0.000 983.920 4.000 ;
    END
  END last_addr[5]
  PIN last_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 992.320 0.000 992.880 4.000 ;
    END
  END last_addr[6]
  PIN last_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1001.280 0.000 1001.840 4.000 ;
    END
  END last_addr[7]
  PIN last_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1010.240 0.000 1010.800 4.000 ;
    END
  END last_addr[8]
  PIN last_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1019.200 0.000 1019.760 4.000 ;
    END
  END last_addr[9]
  PIN le_hi_act
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1062.880 746.000 1063.440 750.000 ;
    END
  END le_hi_act
  PIN le_lo_act
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1042.720 746.000 1043.280 750.000 ;
    END
  END le_lo_act
  PIN ram_bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 649.600 4.000 650.160 ;
    END
  END ram_bus_in[0]
  PIN ram_bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 656.320 4.000 656.880 ;
    END
  END ram_bus_in[1]
  PIN ram_bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 663.040 4.000 663.600 ;
    END
  END ram_bus_in[2]
  PIN ram_bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 669.760 4.000 670.320 ;
    END
  END ram_bus_in[3]
  PIN ram_bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 676.480 4.000 677.040 ;
    END
  END ram_bus_in[4]
  PIN ram_bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 683.200 4.000 683.760 ;
    END
  END ram_bus_in[5]
  PIN ram_bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 689.920 4.000 690.480 ;
    END
  END ram_bus_in[6]
  PIN ram_bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 696.640 4.000 697.200 ;
    END
  END ram_bus_in[7]
  PIN ram_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 703.360 4.000 703.920 ;
    END
  END ram_enabled
  PIN requested_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 619.360 1100.000 619.920 ;
    END
  END requested_addr[0]
  PIN requested_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 686.560 1100.000 687.120 ;
    END
  END requested_addr[10]
  PIN requested_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 693.280 1100.000 693.840 ;
    END
  END requested_addr[11]
  PIN requested_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 700.000 1100.000 700.560 ;
    END
  END requested_addr[12]
  PIN requested_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 706.720 1100.000 707.280 ;
    END
  END requested_addr[13]
  PIN requested_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 713.440 1100.000 714.000 ;
    END
  END requested_addr[14]
  PIN requested_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 720.160 1100.000 720.720 ;
    END
  END requested_addr[15]
  PIN requested_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 626.080 1100.000 626.640 ;
    END
  END requested_addr[1]
  PIN requested_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 632.800 1100.000 633.360 ;
    END
  END requested_addr[2]
  PIN requested_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 639.520 1100.000 640.080 ;
    END
  END requested_addr[3]
  PIN requested_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 646.240 1100.000 646.800 ;
    END
  END requested_addr[4]
  PIN requested_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 652.960 1100.000 653.520 ;
    END
  END requested_addr[5]
  PIN requested_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 659.680 1100.000 660.240 ;
    END
  END requested_addr[6]
  PIN requested_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 666.400 1100.000 666.960 ;
    END
  END requested_addr[7]
  PIN requested_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 673.120 1100.000 673.680 ;
    END
  END requested_addr[8]
  PIN requested_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 679.840 1100.000 680.400 ;
    END
  END requested_addr[9]
  PIN reset_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 484.960 1100.000 485.520 ;
    END
  END reset_out
  PIN rom_bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 595.840 4.000 596.400 ;
    END
  END rom_bus_in[0]
  PIN rom_bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 602.560 4.000 603.120 ;
    END
  END rom_bus_in[1]
  PIN rom_bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 609.280 4.000 609.840 ;
    END
  END rom_bus_in[2]
  PIN rom_bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 616.000 4.000 616.560 ;
    END
  END rom_bus_in[3]
  PIN rom_bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 622.720 4.000 623.280 ;
    END
  END rom_bus_in[4]
  PIN rom_bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 629.440 4.000 630.000 ;
    END
  END rom_bus_in[5]
  PIN rom_bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 636.160 4.000 636.720 ;
    END
  END rom_bus_in[6]
  PIN rom_bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 642.880 4.000 643.440 ;
    END
  END rom_bus_in[7]
  PIN rom_bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 542.080 4.000 542.640 ;
    END
  END rom_bus_out[0]
  PIN rom_bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.800 4.000 549.360 ;
    END
  END rom_bus_out[1]
  PIN rom_bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 555.520 4.000 556.080 ;
    END
  END rom_bus_out[2]
  PIN rom_bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 562.240 4.000 562.800 ;
    END
  END rom_bus_out[3]
  PIN rom_bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 568.960 4.000 569.520 ;
    END
  END rom_bus_out[4]
  PIN rom_bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 575.680 4.000 576.240 ;
    END
  END rom_bus_out[5]
  PIN rom_bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 582.400 4.000 582.960 ;
    END
  END rom_bus_out[6]
  PIN rom_bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 589.120 4.000 589.680 ;
    END
  END rom_bus_out[7]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 733.340 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 733.340 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 0.000 25.200 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 0.000 43.120 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 0.000 374.640 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 0.000 428.400 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 0.000 455.280 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 0.000 509.040 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 0.000 535.920 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 562.240 0.000 562.800 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 589.120 0.000 589.680 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 616.000 0.000 616.560 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 642.880 0.000 643.440 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 0.000 670.320 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 0.000 697.200 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 723.520 0.000 724.080 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 750.400 0.000 750.960 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 777.280 0.000 777.840 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 804.160 0.000 804.720 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 831.040 0.000 831.600 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 857.920 0.000 858.480 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 0.000 132.720 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 884.800 0.000 885.360 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 911.680 0.000 912.240 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 0.000 186.480 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 0.000 213.360 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 0.000 240.240 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 0.000 267.120 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 0.000 294.000 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 0.000 356.720 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 0.000 383.600 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 0.000 410.480 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 0.000 437.360 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 0.000 464.240 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 0.000 491.120 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 0.000 518.000 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 0.000 544.880 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 0.000 571.760 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 0.000 598.640 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 0.000 625.520 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 0.000 652.400 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 0.000 706.160 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 0.000 733.040 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 0.000 759.920 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 0.000 786.800 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 0.000 813.680 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 0.000 840.560 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 0.000 867.440 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 893.760 0.000 894.320 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 920.640 0.000 921.200 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 0.000 222.320 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 0.000 249.200 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 0.000 276.080 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 0.000 302.960 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 0.000 329.840 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 0.000 365.680 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 0.000 392.560 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 0.000 446.320 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 0.000 473.200 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 0.000 500.080 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 0.000 526.960 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 553.280 0.000 553.840 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 0.000 580.720 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 607.040 0.000 607.600 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 0.000 634.480 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 0.000 661.360 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 0.000 688.240 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 0.000 715.120 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 0.000 742.000 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 768.320 0.000 768.880 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 795.200 0.000 795.760 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 0.000 822.640 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 848.960 0.000 849.520 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 875.840 0.000 876.400 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 0.000 150.640 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 902.720 0.000 903.280 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 929.600 0.000 930.160 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 0.000 204.400 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 0.000 231.280 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 0.000 311.920 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 0.000 338.800 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1093.120 734.570 ;
      LAYER Metal2 ;
        RECT 6.860 745.700 34.420 746.000 ;
        RECT 35.580 745.700 54.580 746.000 ;
        RECT 55.740 745.700 74.740 746.000 ;
        RECT 75.900 745.700 94.900 746.000 ;
        RECT 96.060 745.700 115.060 746.000 ;
        RECT 116.220 745.700 135.220 746.000 ;
        RECT 136.380 745.700 155.380 746.000 ;
        RECT 156.540 745.700 175.540 746.000 ;
        RECT 176.700 745.700 195.700 746.000 ;
        RECT 196.860 745.700 215.860 746.000 ;
        RECT 217.020 745.700 236.020 746.000 ;
        RECT 237.180 745.700 256.180 746.000 ;
        RECT 257.340 745.700 276.340 746.000 ;
        RECT 277.500 745.700 296.500 746.000 ;
        RECT 297.660 745.700 316.660 746.000 ;
        RECT 317.820 745.700 336.820 746.000 ;
        RECT 337.980 745.700 356.980 746.000 ;
        RECT 358.140 745.700 377.140 746.000 ;
        RECT 378.300 745.700 397.300 746.000 ;
        RECT 398.460 745.700 417.460 746.000 ;
        RECT 418.620 745.700 437.620 746.000 ;
        RECT 438.780 745.700 457.780 746.000 ;
        RECT 458.940 745.700 477.940 746.000 ;
        RECT 479.100 745.700 498.100 746.000 ;
        RECT 499.260 745.700 518.260 746.000 ;
        RECT 519.420 745.700 538.420 746.000 ;
        RECT 539.580 745.700 558.580 746.000 ;
        RECT 559.740 745.700 578.740 746.000 ;
        RECT 579.900 745.700 598.900 746.000 ;
        RECT 600.060 745.700 619.060 746.000 ;
        RECT 620.220 745.700 639.220 746.000 ;
        RECT 640.380 745.700 659.380 746.000 ;
        RECT 660.540 745.700 679.540 746.000 ;
        RECT 680.700 745.700 699.700 746.000 ;
        RECT 700.860 745.700 719.860 746.000 ;
        RECT 721.020 745.700 740.020 746.000 ;
        RECT 741.180 745.700 760.180 746.000 ;
        RECT 761.340 745.700 780.340 746.000 ;
        RECT 781.500 745.700 800.500 746.000 ;
        RECT 801.660 745.700 820.660 746.000 ;
        RECT 821.820 745.700 840.820 746.000 ;
        RECT 841.980 745.700 860.980 746.000 ;
        RECT 862.140 745.700 881.140 746.000 ;
        RECT 882.300 745.700 901.300 746.000 ;
        RECT 902.460 745.700 921.460 746.000 ;
        RECT 922.620 745.700 941.620 746.000 ;
        RECT 942.780 745.700 961.780 746.000 ;
        RECT 962.940 745.700 981.940 746.000 ;
        RECT 983.100 745.700 1002.100 746.000 ;
        RECT 1003.260 745.700 1022.260 746.000 ;
        RECT 1023.420 745.700 1042.420 746.000 ;
        RECT 1043.580 745.700 1062.580 746.000 ;
        RECT 1063.740 745.700 1091.860 746.000 ;
        RECT 6.860 4.300 1091.860 745.700 ;
        RECT 6.860 3.500 24.340 4.300 ;
        RECT 25.500 3.500 33.300 4.300 ;
        RECT 34.460 3.500 42.260 4.300 ;
        RECT 43.420 3.500 51.220 4.300 ;
        RECT 52.380 3.500 60.180 4.300 ;
        RECT 61.340 3.500 69.140 4.300 ;
        RECT 70.300 3.500 78.100 4.300 ;
        RECT 79.260 3.500 87.060 4.300 ;
        RECT 88.220 3.500 96.020 4.300 ;
        RECT 97.180 3.500 104.980 4.300 ;
        RECT 106.140 3.500 113.940 4.300 ;
        RECT 115.100 3.500 122.900 4.300 ;
        RECT 124.060 3.500 131.860 4.300 ;
        RECT 133.020 3.500 140.820 4.300 ;
        RECT 141.980 3.500 149.780 4.300 ;
        RECT 150.940 3.500 158.740 4.300 ;
        RECT 159.900 3.500 167.700 4.300 ;
        RECT 168.860 3.500 176.660 4.300 ;
        RECT 177.820 3.500 185.620 4.300 ;
        RECT 186.780 3.500 194.580 4.300 ;
        RECT 195.740 3.500 203.540 4.300 ;
        RECT 204.700 3.500 212.500 4.300 ;
        RECT 213.660 3.500 221.460 4.300 ;
        RECT 222.620 3.500 230.420 4.300 ;
        RECT 231.580 3.500 239.380 4.300 ;
        RECT 240.540 3.500 248.340 4.300 ;
        RECT 249.500 3.500 257.300 4.300 ;
        RECT 258.460 3.500 266.260 4.300 ;
        RECT 267.420 3.500 275.220 4.300 ;
        RECT 276.380 3.500 284.180 4.300 ;
        RECT 285.340 3.500 293.140 4.300 ;
        RECT 294.300 3.500 302.100 4.300 ;
        RECT 303.260 3.500 311.060 4.300 ;
        RECT 312.220 3.500 320.020 4.300 ;
        RECT 321.180 3.500 328.980 4.300 ;
        RECT 330.140 3.500 337.940 4.300 ;
        RECT 339.100 3.500 346.900 4.300 ;
        RECT 348.060 3.500 355.860 4.300 ;
        RECT 357.020 3.500 364.820 4.300 ;
        RECT 365.980 3.500 373.780 4.300 ;
        RECT 374.940 3.500 382.740 4.300 ;
        RECT 383.900 3.500 391.700 4.300 ;
        RECT 392.860 3.500 400.660 4.300 ;
        RECT 401.820 3.500 409.620 4.300 ;
        RECT 410.780 3.500 418.580 4.300 ;
        RECT 419.740 3.500 427.540 4.300 ;
        RECT 428.700 3.500 436.500 4.300 ;
        RECT 437.660 3.500 445.460 4.300 ;
        RECT 446.620 3.500 454.420 4.300 ;
        RECT 455.580 3.500 463.380 4.300 ;
        RECT 464.540 3.500 472.340 4.300 ;
        RECT 473.500 3.500 481.300 4.300 ;
        RECT 482.460 3.500 490.260 4.300 ;
        RECT 491.420 3.500 499.220 4.300 ;
        RECT 500.380 3.500 508.180 4.300 ;
        RECT 509.340 3.500 517.140 4.300 ;
        RECT 518.300 3.500 526.100 4.300 ;
        RECT 527.260 3.500 535.060 4.300 ;
        RECT 536.220 3.500 544.020 4.300 ;
        RECT 545.180 3.500 552.980 4.300 ;
        RECT 554.140 3.500 561.940 4.300 ;
        RECT 563.100 3.500 570.900 4.300 ;
        RECT 572.060 3.500 579.860 4.300 ;
        RECT 581.020 3.500 588.820 4.300 ;
        RECT 589.980 3.500 597.780 4.300 ;
        RECT 598.940 3.500 606.740 4.300 ;
        RECT 607.900 3.500 615.700 4.300 ;
        RECT 616.860 3.500 624.660 4.300 ;
        RECT 625.820 3.500 633.620 4.300 ;
        RECT 634.780 3.500 642.580 4.300 ;
        RECT 643.740 3.500 651.540 4.300 ;
        RECT 652.700 3.500 660.500 4.300 ;
        RECT 661.660 3.500 669.460 4.300 ;
        RECT 670.620 3.500 678.420 4.300 ;
        RECT 679.580 3.500 687.380 4.300 ;
        RECT 688.540 3.500 696.340 4.300 ;
        RECT 697.500 3.500 705.300 4.300 ;
        RECT 706.460 3.500 714.260 4.300 ;
        RECT 715.420 3.500 723.220 4.300 ;
        RECT 724.380 3.500 732.180 4.300 ;
        RECT 733.340 3.500 741.140 4.300 ;
        RECT 742.300 3.500 750.100 4.300 ;
        RECT 751.260 3.500 759.060 4.300 ;
        RECT 760.220 3.500 768.020 4.300 ;
        RECT 769.180 3.500 776.980 4.300 ;
        RECT 778.140 3.500 785.940 4.300 ;
        RECT 787.100 3.500 794.900 4.300 ;
        RECT 796.060 3.500 803.860 4.300 ;
        RECT 805.020 3.500 812.820 4.300 ;
        RECT 813.980 3.500 821.780 4.300 ;
        RECT 822.940 3.500 830.740 4.300 ;
        RECT 831.900 3.500 839.700 4.300 ;
        RECT 840.860 3.500 848.660 4.300 ;
        RECT 849.820 3.500 857.620 4.300 ;
        RECT 858.780 3.500 866.580 4.300 ;
        RECT 867.740 3.500 875.540 4.300 ;
        RECT 876.700 3.500 884.500 4.300 ;
        RECT 885.660 3.500 893.460 4.300 ;
        RECT 894.620 3.500 902.420 4.300 ;
        RECT 903.580 3.500 911.380 4.300 ;
        RECT 912.540 3.500 920.340 4.300 ;
        RECT 921.500 3.500 929.300 4.300 ;
        RECT 930.460 3.500 938.260 4.300 ;
        RECT 939.420 3.500 947.220 4.300 ;
        RECT 948.380 3.500 956.180 4.300 ;
        RECT 957.340 3.500 965.140 4.300 ;
        RECT 966.300 3.500 974.100 4.300 ;
        RECT 975.260 3.500 983.060 4.300 ;
        RECT 984.220 3.500 992.020 4.300 ;
        RECT 993.180 3.500 1000.980 4.300 ;
        RECT 1002.140 3.500 1009.940 4.300 ;
        RECT 1011.100 3.500 1018.900 4.300 ;
        RECT 1020.060 3.500 1027.860 4.300 ;
        RECT 1029.020 3.500 1036.820 4.300 ;
        RECT 1037.980 3.500 1045.780 4.300 ;
        RECT 1046.940 3.500 1054.740 4.300 ;
        RECT 1055.900 3.500 1063.700 4.300 ;
        RECT 1064.860 3.500 1072.660 4.300 ;
        RECT 1073.820 3.500 1091.860 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 721.020 1096.340 733.180 ;
        RECT 4.000 719.860 1095.700 721.020 ;
        RECT 4.000 714.300 1096.340 719.860 ;
        RECT 4.000 713.140 1095.700 714.300 ;
        RECT 4.000 707.580 1096.340 713.140 ;
        RECT 4.000 706.420 1095.700 707.580 ;
        RECT 4.000 704.220 1096.340 706.420 ;
        RECT 4.300 703.060 1096.340 704.220 ;
        RECT 4.000 700.860 1096.340 703.060 ;
        RECT 4.000 699.700 1095.700 700.860 ;
        RECT 4.000 697.500 1096.340 699.700 ;
        RECT 4.300 696.340 1096.340 697.500 ;
        RECT 4.000 694.140 1096.340 696.340 ;
        RECT 4.000 692.980 1095.700 694.140 ;
        RECT 4.000 690.780 1096.340 692.980 ;
        RECT 4.300 689.620 1096.340 690.780 ;
        RECT 4.000 687.420 1096.340 689.620 ;
        RECT 4.000 686.260 1095.700 687.420 ;
        RECT 4.000 684.060 1096.340 686.260 ;
        RECT 4.300 682.900 1096.340 684.060 ;
        RECT 4.000 680.700 1096.340 682.900 ;
        RECT 4.000 679.540 1095.700 680.700 ;
        RECT 4.000 677.340 1096.340 679.540 ;
        RECT 4.300 676.180 1096.340 677.340 ;
        RECT 4.000 673.980 1096.340 676.180 ;
        RECT 4.000 672.820 1095.700 673.980 ;
        RECT 4.000 670.620 1096.340 672.820 ;
        RECT 4.300 669.460 1096.340 670.620 ;
        RECT 4.000 667.260 1096.340 669.460 ;
        RECT 4.000 666.100 1095.700 667.260 ;
        RECT 4.000 663.900 1096.340 666.100 ;
        RECT 4.300 662.740 1096.340 663.900 ;
        RECT 4.000 660.540 1096.340 662.740 ;
        RECT 4.000 659.380 1095.700 660.540 ;
        RECT 4.000 657.180 1096.340 659.380 ;
        RECT 4.300 656.020 1096.340 657.180 ;
        RECT 4.000 653.820 1096.340 656.020 ;
        RECT 4.000 652.660 1095.700 653.820 ;
        RECT 4.000 650.460 1096.340 652.660 ;
        RECT 4.300 649.300 1096.340 650.460 ;
        RECT 4.000 647.100 1096.340 649.300 ;
        RECT 4.000 645.940 1095.700 647.100 ;
        RECT 4.000 643.740 1096.340 645.940 ;
        RECT 4.300 642.580 1096.340 643.740 ;
        RECT 4.000 640.380 1096.340 642.580 ;
        RECT 4.000 639.220 1095.700 640.380 ;
        RECT 4.000 637.020 1096.340 639.220 ;
        RECT 4.300 635.860 1096.340 637.020 ;
        RECT 4.000 633.660 1096.340 635.860 ;
        RECT 4.000 632.500 1095.700 633.660 ;
        RECT 4.000 630.300 1096.340 632.500 ;
        RECT 4.300 629.140 1096.340 630.300 ;
        RECT 4.000 626.940 1096.340 629.140 ;
        RECT 4.000 625.780 1095.700 626.940 ;
        RECT 4.000 623.580 1096.340 625.780 ;
        RECT 4.300 622.420 1096.340 623.580 ;
        RECT 4.000 620.220 1096.340 622.420 ;
        RECT 4.000 619.060 1095.700 620.220 ;
        RECT 4.000 616.860 1096.340 619.060 ;
        RECT 4.300 615.700 1096.340 616.860 ;
        RECT 4.000 613.500 1096.340 615.700 ;
        RECT 4.000 612.340 1095.700 613.500 ;
        RECT 4.000 610.140 1096.340 612.340 ;
        RECT 4.300 608.980 1096.340 610.140 ;
        RECT 4.000 606.780 1096.340 608.980 ;
        RECT 4.000 605.620 1095.700 606.780 ;
        RECT 4.000 603.420 1096.340 605.620 ;
        RECT 4.300 602.260 1096.340 603.420 ;
        RECT 4.000 600.060 1096.340 602.260 ;
        RECT 4.000 598.900 1095.700 600.060 ;
        RECT 4.000 596.700 1096.340 598.900 ;
        RECT 4.300 595.540 1096.340 596.700 ;
        RECT 4.000 593.340 1096.340 595.540 ;
        RECT 4.000 592.180 1095.700 593.340 ;
        RECT 4.000 589.980 1096.340 592.180 ;
        RECT 4.300 588.820 1096.340 589.980 ;
        RECT 4.000 586.620 1096.340 588.820 ;
        RECT 4.000 585.460 1095.700 586.620 ;
        RECT 4.000 583.260 1096.340 585.460 ;
        RECT 4.300 582.100 1096.340 583.260 ;
        RECT 4.000 579.900 1096.340 582.100 ;
        RECT 4.000 578.740 1095.700 579.900 ;
        RECT 4.000 576.540 1096.340 578.740 ;
        RECT 4.300 575.380 1096.340 576.540 ;
        RECT 4.000 573.180 1096.340 575.380 ;
        RECT 4.000 572.020 1095.700 573.180 ;
        RECT 4.000 569.820 1096.340 572.020 ;
        RECT 4.300 568.660 1096.340 569.820 ;
        RECT 4.000 566.460 1096.340 568.660 ;
        RECT 4.000 565.300 1095.700 566.460 ;
        RECT 4.000 563.100 1096.340 565.300 ;
        RECT 4.300 561.940 1096.340 563.100 ;
        RECT 4.000 559.740 1096.340 561.940 ;
        RECT 4.000 558.580 1095.700 559.740 ;
        RECT 4.000 556.380 1096.340 558.580 ;
        RECT 4.300 555.220 1096.340 556.380 ;
        RECT 4.000 553.020 1096.340 555.220 ;
        RECT 4.000 551.860 1095.700 553.020 ;
        RECT 4.000 549.660 1096.340 551.860 ;
        RECT 4.300 548.500 1096.340 549.660 ;
        RECT 4.000 546.300 1096.340 548.500 ;
        RECT 4.000 545.140 1095.700 546.300 ;
        RECT 4.000 542.940 1096.340 545.140 ;
        RECT 4.300 541.780 1096.340 542.940 ;
        RECT 4.000 539.580 1096.340 541.780 ;
        RECT 4.000 538.420 1095.700 539.580 ;
        RECT 4.000 536.220 1096.340 538.420 ;
        RECT 4.300 535.060 1096.340 536.220 ;
        RECT 4.000 532.860 1096.340 535.060 ;
        RECT 4.000 531.700 1095.700 532.860 ;
        RECT 4.000 529.500 1096.340 531.700 ;
        RECT 4.300 528.340 1096.340 529.500 ;
        RECT 4.000 526.140 1096.340 528.340 ;
        RECT 4.000 524.980 1095.700 526.140 ;
        RECT 4.000 522.780 1096.340 524.980 ;
        RECT 4.300 521.620 1096.340 522.780 ;
        RECT 4.000 519.420 1096.340 521.620 ;
        RECT 4.000 518.260 1095.700 519.420 ;
        RECT 4.000 516.060 1096.340 518.260 ;
        RECT 4.300 514.900 1096.340 516.060 ;
        RECT 4.000 512.700 1096.340 514.900 ;
        RECT 4.000 511.540 1095.700 512.700 ;
        RECT 4.000 509.340 1096.340 511.540 ;
        RECT 4.300 508.180 1096.340 509.340 ;
        RECT 4.000 505.980 1096.340 508.180 ;
        RECT 4.000 504.820 1095.700 505.980 ;
        RECT 4.000 502.620 1096.340 504.820 ;
        RECT 4.300 501.460 1096.340 502.620 ;
        RECT 4.000 499.260 1096.340 501.460 ;
        RECT 4.000 498.100 1095.700 499.260 ;
        RECT 4.000 495.900 1096.340 498.100 ;
        RECT 4.300 494.740 1096.340 495.900 ;
        RECT 4.000 492.540 1096.340 494.740 ;
        RECT 4.000 491.380 1095.700 492.540 ;
        RECT 4.000 489.180 1096.340 491.380 ;
        RECT 4.300 488.020 1096.340 489.180 ;
        RECT 4.000 485.820 1096.340 488.020 ;
        RECT 4.000 484.660 1095.700 485.820 ;
        RECT 4.000 482.460 1096.340 484.660 ;
        RECT 4.300 481.300 1096.340 482.460 ;
        RECT 4.000 479.100 1096.340 481.300 ;
        RECT 4.000 477.940 1095.700 479.100 ;
        RECT 4.000 475.740 1096.340 477.940 ;
        RECT 4.300 474.580 1096.340 475.740 ;
        RECT 4.000 472.380 1096.340 474.580 ;
        RECT 4.000 471.220 1095.700 472.380 ;
        RECT 4.000 469.020 1096.340 471.220 ;
        RECT 4.300 467.860 1096.340 469.020 ;
        RECT 4.000 465.660 1096.340 467.860 ;
        RECT 4.000 464.500 1095.700 465.660 ;
        RECT 4.000 462.300 1096.340 464.500 ;
        RECT 4.300 461.140 1096.340 462.300 ;
        RECT 4.000 458.940 1096.340 461.140 ;
        RECT 4.000 457.780 1095.700 458.940 ;
        RECT 4.000 455.580 1096.340 457.780 ;
        RECT 4.300 454.420 1096.340 455.580 ;
        RECT 4.000 452.220 1096.340 454.420 ;
        RECT 4.000 451.060 1095.700 452.220 ;
        RECT 4.000 448.860 1096.340 451.060 ;
        RECT 4.300 447.700 1096.340 448.860 ;
        RECT 4.000 445.500 1096.340 447.700 ;
        RECT 4.000 444.340 1095.700 445.500 ;
        RECT 4.000 442.140 1096.340 444.340 ;
        RECT 4.300 440.980 1096.340 442.140 ;
        RECT 4.000 438.780 1096.340 440.980 ;
        RECT 4.000 437.620 1095.700 438.780 ;
        RECT 4.000 435.420 1096.340 437.620 ;
        RECT 4.300 434.260 1096.340 435.420 ;
        RECT 4.000 432.060 1096.340 434.260 ;
        RECT 4.000 430.900 1095.700 432.060 ;
        RECT 4.000 428.700 1096.340 430.900 ;
        RECT 4.300 427.540 1096.340 428.700 ;
        RECT 4.000 425.340 1096.340 427.540 ;
        RECT 4.000 424.180 1095.700 425.340 ;
        RECT 4.000 421.980 1096.340 424.180 ;
        RECT 4.300 420.820 1096.340 421.980 ;
        RECT 4.000 418.620 1096.340 420.820 ;
        RECT 4.000 417.460 1095.700 418.620 ;
        RECT 4.000 415.260 1096.340 417.460 ;
        RECT 4.300 414.100 1096.340 415.260 ;
        RECT 4.000 411.900 1096.340 414.100 ;
        RECT 4.000 410.740 1095.700 411.900 ;
        RECT 4.000 408.540 1096.340 410.740 ;
        RECT 4.300 407.380 1096.340 408.540 ;
        RECT 4.000 405.180 1096.340 407.380 ;
        RECT 4.000 404.020 1095.700 405.180 ;
        RECT 4.000 401.820 1096.340 404.020 ;
        RECT 4.300 400.660 1096.340 401.820 ;
        RECT 4.000 398.460 1096.340 400.660 ;
        RECT 4.000 397.300 1095.700 398.460 ;
        RECT 4.000 395.100 1096.340 397.300 ;
        RECT 4.300 393.940 1096.340 395.100 ;
        RECT 4.000 391.740 1096.340 393.940 ;
        RECT 4.000 390.580 1095.700 391.740 ;
        RECT 4.000 388.380 1096.340 390.580 ;
        RECT 4.300 387.220 1096.340 388.380 ;
        RECT 4.000 385.020 1096.340 387.220 ;
        RECT 4.000 383.860 1095.700 385.020 ;
        RECT 4.000 381.660 1096.340 383.860 ;
        RECT 4.300 380.500 1096.340 381.660 ;
        RECT 4.000 378.300 1096.340 380.500 ;
        RECT 4.000 377.140 1095.700 378.300 ;
        RECT 4.000 374.940 1096.340 377.140 ;
        RECT 4.300 373.780 1096.340 374.940 ;
        RECT 4.000 371.580 1096.340 373.780 ;
        RECT 4.000 370.420 1095.700 371.580 ;
        RECT 4.000 368.220 1096.340 370.420 ;
        RECT 4.300 367.060 1096.340 368.220 ;
        RECT 4.000 364.860 1096.340 367.060 ;
        RECT 4.000 363.700 1095.700 364.860 ;
        RECT 4.000 361.500 1096.340 363.700 ;
        RECT 4.300 360.340 1096.340 361.500 ;
        RECT 4.000 358.140 1096.340 360.340 ;
        RECT 4.000 356.980 1095.700 358.140 ;
        RECT 4.000 354.780 1096.340 356.980 ;
        RECT 4.300 353.620 1096.340 354.780 ;
        RECT 4.000 351.420 1096.340 353.620 ;
        RECT 4.000 350.260 1095.700 351.420 ;
        RECT 4.000 348.060 1096.340 350.260 ;
        RECT 4.300 346.900 1096.340 348.060 ;
        RECT 4.000 344.700 1096.340 346.900 ;
        RECT 4.000 343.540 1095.700 344.700 ;
        RECT 4.000 341.340 1096.340 343.540 ;
        RECT 4.300 340.180 1096.340 341.340 ;
        RECT 4.000 337.980 1096.340 340.180 ;
        RECT 4.000 336.820 1095.700 337.980 ;
        RECT 4.000 334.620 1096.340 336.820 ;
        RECT 4.300 333.460 1096.340 334.620 ;
        RECT 4.000 331.260 1096.340 333.460 ;
        RECT 4.000 330.100 1095.700 331.260 ;
        RECT 4.000 327.900 1096.340 330.100 ;
        RECT 4.300 326.740 1096.340 327.900 ;
        RECT 4.000 324.540 1096.340 326.740 ;
        RECT 4.000 323.380 1095.700 324.540 ;
        RECT 4.000 321.180 1096.340 323.380 ;
        RECT 4.300 320.020 1096.340 321.180 ;
        RECT 4.000 317.820 1096.340 320.020 ;
        RECT 4.000 316.660 1095.700 317.820 ;
        RECT 4.000 314.460 1096.340 316.660 ;
        RECT 4.300 313.300 1096.340 314.460 ;
        RECT 4.000 311.100 1096.340 313.300 ;
        RECT 4.000 309.940 1095.700 311.100 ;
        RECT 4.000 307.740 1096.340 309.940 ;
        RECT 4.300 306.580 1096.340 307.740 ;
        RECT 4.000 304.380 1096.340 306.580 ;
        RECT 4.000 303.220 1095.700 304.380 ;
        RECT 4.000 301.020 1096.340 303.220 ;
        RECT 4.300 299.860 1096.340 301.020 ;
        RECT 4.000 297.660 1096.340 299.860 ;
        RECT 4.000 296.500 1095.700 297.660 ;
        RECT 4.000 294.300 1096.340 296.500 ;
        RECT 4.300 293.140 1096.340 294.300 ;
        RECT 4.000 290.940 1096.340 293.140 ;
        RECT 4.000 289.780 1095.700 290.940 ;
        RECT 4.000 287.580 1096.340 289.780 ;
        RECT 4.300 286.420 1096.340 287.580 ;
        RECT 4.000 284.220 1096.340 286.420 ;
        RECT 4.000 283.060 1095.700 284.220 ;
        RECT 4.000 280.860 1096.340 283.060 ;
        RECT 4.300 279.700 1096.340 280.860 ;
        RECT 4.000 277.500 1096.340 279.700 ;
        RECT 4.000 276.340 1095.700 277.500 ;
        RECT 4.000 274.140 1096.340 276.340 ;
        RECT 4.300 272.980 1096.340 274.140 ;
        RECT 4.000 270.780 1096.340 272.980 ;
        RECT 4.000 269.620 1095.700 270.780 ;
        RECT 4.000 267.420 1096.340 269.620 ;
        RECT 4.300 266.260 1096.340 267.420 ;
        RECT 4.000 264.060 1096.340 266.260 ;
        RECT 4.000 262.900 1095.700 264.060 ;
        RECT 4.000 260.700 1096.340 262.900 ;
        RECT 4.300 259.540 1096.340 260.700 ;
        RECT 4.000 257.340 1096.340 259.540 ;
        RECT 4.000 256.180 1095.700 257.340 ;
        RECT 4.000 253.980 1096.340 256.180 ;
        RECT 4.300 252.820 1096.340 253.980 ;
        RECT 4.000 250.620 1096.340 252.820 ;
        RECT 4.000 249.460 1095.700 250.620 ;
        RECT 4.000 247.260 1096.340 249.460 ;
        RECT 4.300 246.100 1096.340 247.260 ;
        RECT 4.000 243.900 1096.340 246.100 ;
        RECT 4.000 242.740 1095.700 243.900 ;
        RECT 4.000 240.540 1096.340 242.740 ;
        RECT 4.300 239.380 1096.340 240.540 ;
        RECT 4.000 237.180 1096.340 239.380 ;
        RECT 4.000 236.020 1095.700 237.180 ;
        RECT 4.000 233.820 1096.340 236.020 ;
        RECT 4.300 232.660 1096.340 233.820 ;
        RECT 4.000 230.460 1096.340 232.660 ;
        RECT 4.000 229.300 1095.700 230.460 ;
        RECT 4.000 227.100 1096.340 229.300 ;
        RECT 4.300 225.940 1096.340 227.100 ;
        RECT 4.000 223.740 1096.340 225.940 ;
        RECT 4.000 222.580 1095.700 223.740 ;
        RECT 4.000 220.380 1096.340 222.580 ;
        RECT 4.300 219.220 1096.340 220.380 ;
        RECT 4.000 217.020 1096.340 219.220 ;
        RECT 4.000 215.860 1095.700 217.020 ;
        RECT 4.000 213.660 1096.340 215.860 ;
        RECT 4.300 212.500 1096.340 213.660 ;
        RECT 4.000 210.300 1096.340 212.500 ;
        RECT 4.000 209.140 1095.700 210.300 ;
        RECT 4.000 206.940 1096.340 209.140 ;
        RECT 4.300 205.780 1096.340 206.940 ;
        RECT 4.000 203.580 1096.340 205.780 ;
        RECT 4.000 202.420 1095.700 203.580 ;
        RECT 4.000 200.220 1096.340 202.420 ;
        RECT 4.300 199.060 1096.340 200.220 ;
        RECT 4.000 196.860 1096.340 199.060 ;
        RECT 4.000 195.700 1095.700 196.860 ;
        RECT 4.000 193.500 1096.340 195.700 ;
        RECT 4.300 192.340 1096.340 193.500 ;
        RECT 4.000 190.140 1096.340 192.340 ;
        RECT 4.000 188.980 1095.700 190.140 ;
        RECT 4.000 186.780 1096.340 188.980 ;
        RECT 4.300 185.620 1096.340 186.780 ;
        RECT 4.000 183.420 1096.340 185.620 ;
        RECT 4.000 182.260 1095.700 183.420 ;
        RECT 4.000 180.060 1096.340 182.260 ;
        RECT 4.300 178.900 1096.340 180.060 ;
        RECT 4.000 176.700 1096.340 178.900 ;
        RECT 4.000 175.540 1095.700 176.700 ;
        RECT 4.000 173.340 1096.340 175.540 ;
        RECT 4.300 172.180 1096.340 173.340 ;
        RECT 4.000 169.980 1096.340 172.180 ;
        RECT 4.000 168.820 1095.700 169.980 ;
        RECT 4.000 166.620 1096.340 168.820 ;
        RECT 4.300 165.460 1096.340 166.620 ;
        RECT 4.000 163.260 1096.340 165.460 ;
        RECT 4.000 162.100 1095.700 163.260 ;
        RECT 4.000 159.900 1096.340 162.100 ;
        RECT 4.300 158.740 1096.340 159.900 ;
        RECT 4.000 156.540 1096.340 158.740 ;
        RECT 4.000 155.380 1095.700 156.540 ;
        RECT 4.000 153.180 1096.340 155.380 ;
        RECT 4.300 152.020 1096.340 153.180 ;
        RECT 4.000 149.820 1096.340 152.020 ;
        RECT 4.000 148.660 1095.700 149.820 ;
        RECT 4.000 146.460 1096.340 148.660 ;
        RECT 4.300 145.300 1096.340 146.460 ;
        RECT 4.000 143.100 1096.340 145.300 ;
        RECT 4.000 141.940 1095.700 143.100 ;
        RECT 4.000 139.740 1096.340 141.940 ;
        RECT 4.300 138.580 1096.340 139.740 ;
        RECT 4.000 136.380 1096.340 138.580 ;
        RECT 4.000 135.220 1095.700 136.380 ;
        RECT 4.000 133.020 1096.340 135.220 ;
        RECT 4.300 131.860 1096.340 133.020 ;
        RECT 4.000 129.660 1096.340 131.860 ;
        RECT 4.000 128.500 1095.700 129.660 ;
        RECT 4.000 126.300 1096.340 128.500 ;
        RECT 4.300 125.140 1096.340 126.300 ;
        RECT 4.000 122.940 1096.340 125.140 ;
        RECT 4.000 121.780 1095.700 122.940 ;
        RECT 4.000 119.580 1096.340 121.780 ;
        RECT 4.300 118.420 1096.340 119.580 ;
        RECT 4.000 116.220 1096.340 118.420 ;
        RECT 4.000 115.060 1095.700 116.220 ;
        RECT 4.000 112.860 1096.340 115.060 ;
        RECT 4.300 111.700 1096.340 112.860 ;
        RECT 4.000 109.500 1096.340 111.700 ;
        RECT 4.000 108.340 1095.700 109.500 ;
        RECT 4.000 106.140 1096.340 108.340 ;
        RECT 4.300 104.980 1096.340 106.140 ;
        RECT 4.000 102.780 1096.340 104.980 ;
        RECT 4.000 101.620 1095.700 102.780 ;
        RECT 4.000 99.420 1096.340 101.620 ;
        RECT 4.300 98.260 1096.340 99.420 ;
        RECT 4.000 96.060 1096.340 98.260 ;
        RECT 4.000 94.900 1095.700 96.060 ;
        RECT 4.000 92.700 1096.340 94.900 ;
        RECT 4.300 91.540 1096.340 92.700 ;
        RECT 4.000 89.340 1096.340 91.540 ;
        RECT 4.000 88.180 1095.700 89.340 ;
        RECT 4.000 85.980 1096.340 88.180 ;
        RECT 4.300 84.820 1096.340 85.980 ;
        RECT 4.000 82.620 1096.340 84.820 ;
        RECT 4.000 81.460 1095.700 82.620 ;
        RECT 4.000 79.260 1096.340 81.460 ;
        RECT 4.300 78.100 1096.340 79.260 ;
        RECT 4.000 75.900 1096.340 78.100 ;
        RECT 4.000 74.740 1095.700 75.900 ;
        RECT 4.000 72.540 1096.340 74.740 ;
        RECT 4.300 71.380 1096.340 72.540 ;
        RECT 4.000 69.180 1096.340 71.380 ;
        RECT 4.000 68.020 1095.700 69.180 ;
        RECT 4.000 65.820 1096.340 68.020 ;
        RECT 4.300 64.660 1096.340 65.820 ;
        RECT 4.000 62.460 1096.340 64.660 ;
        RECT 4.000 61.300 1095.700 62.460 ;
        RECT 4.000 59.100 1096.340 61.300 ;
        RECT 4.300 57.940 1096.340 59.100 ;
        RECT 4.000 55.740 1096.340 57.940 ;
        RECT 4.000 54.580 1095.700 55.740 ;
        RECT 4.000 52.380 1096.340 54.580 ;
        RECT 4.300 51.220 1096.340 52.380 ;
        RECT 4.000 49.020 1096.340 51.220 ;
        RECT 4.000 47.860 1095.700 49.020 ;
        RECT 4.000 45.660 1096.340 47.860 ;
        RECT 4.300 44.500 1096.340 45.660 ;
        RECT 4.000 42.300 1096.340 44.500 ;
        RECT 4.000 41.140 1095.700 42.300 ;
        RECT 4.000 35.580 1096.340 41.140 ;
        RECT 4.000 34.420 1095.700 35.580 ;
        RECT 4.000 28.860 1096.340 34.420 ;
        RECT 4.000 27.700 1095.700 28.860 ;
        RECT 4.000 13.580 1096.340 27.700 ;
      LAYER Metal4 ;
        RECT 18.620 17.450 21.940 640.550 ;
        RECT 24.140 17.450 98.740 640.550 ;
        RECT 100.940 17.450 175.540 640.550 ;
        RECT 177.740 17.450 252.340 640.550 ;
        RECT 254.540 17.450 329.140 640.550 ;
        RECT 331.340 17.450 405.940 640.550 ;
        RECT 408.140 17.450 482.740 640.550 ;
        RECT 484.940 17.450 559.540 640.550 ;
        RECT 561.740 17.450 636.340 640.550 ;
        RECT 638.540 17.450 713.140 640.550 ;
        RECT 715.340 17.450 789.940 640.550 ;
        RECT 792.140 17.450 866.740 640.550 ;
        RECT 868.940 17.450 943.540 640.550 ;
        RECT 945.740 17.450 1020.340 640.550 ;
        RECT 1022.540 17.450 1081.780 640.550 ;
  END
END wrapped_as2650
END LIBRARY

