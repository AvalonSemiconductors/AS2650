VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as2650
  CLASS BLOCK ;
  FOREIGN wrapped_as2650 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 800.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 796.000 43.120 800.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 796.000 311.920 800.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 796.000 338.800 800.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 796.000 365.680 800.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 796.000 392.560 800.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 796.000 419.440 800.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 796.000 446.320 800.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 796.000 473.200 800.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 796.000 500.080 800.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 796.000 526.960 800.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 553.280 796.000 553.840 800.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 796.000 70.000 800.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 796.000 580.720 800.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 607.040 796.000 607.600 800.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 796.000 634.480 800.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 796.000 661.360 800.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 796.000 688.240 800.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 796.000 715.120 800.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 796.000 742.000 800.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 768.320 796.000 768.880 800.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 795.200 796.000 795.760 800.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 796.000 822.640 800.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 796.000 96.880 800.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 848.960 796.000 849.520 800.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 875.840 796.000 876.400 800.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 902.720 796.000 903.280 800.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 929.600 796.000 930.160 800.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 956.480 796.000 957.040 800.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 796.000 983.920 800.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1010.240 796.000 1010.800 800.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1037.120 796.000 1037.680 800.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 796.000 123.760 800.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 796.000 150.640 800.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 796.000 177.520 800.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 796.000 204.400 800.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 796.000 231.280 800.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 796.000 258.160 800.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 796.000 285.040 800.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 796.000 52.080 800.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 796.000 320.880 800.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 796.000 347.760 800.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 796.000 374.640 800.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 796.000 401.520 800.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 796.000 428.400 800.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 796.000 455.280 800.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 796.000 482.160 800.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 796.000 509.040 800.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 796.000 535.920 800.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 562.240 796.000 562.800 800.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 796.000 78.960 800.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 589.120 796.000 589.680 800.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 616.000 796.000 616.560 800.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 642.880 796.000 643.440 800.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 796.000 670.320 800.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 796.000 697.200 800.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 723.520 796.000 724.080 800.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 750.400 796.000 750.960 800.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 777.280 796.000 777.840 800.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 804.160 796.000 804.720 800.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 831.040 796.000 831.600 800.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 796.000 105.840 800.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 857.920 796.000 858.480 800.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 884.800 796.000 885.360 800.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 911.680 796.000 912.240 800.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 938.560 796.000 939.120 800.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 965.440 796.000 966.000 800.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 992.320 796.000 992.880 800.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1019.200 796.000 1019.760 800.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1046.080 796.000 1046.640 800.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 796.000 132.720 800.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 796.000 159.600 800.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 796.000 186.480 800.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 796.000 213.360 800.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 796.000 240.240 800.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 796.000 267.120 800.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 796.000 294.000 800.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 796.000 61.040 800.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 796.000 329.840 800.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 796.000 356.720 800.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 796.000 383.600 800.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 796.000 410.480 800.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 796.000 437.360 800.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 796.000 464.240 800.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 796.000 491.120 800.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 796.000 518.000 800.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 796.000 544.880 800.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 796.000 571.760 800.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 796.000 87.920 800.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 796.000 598.640 800.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 796.000 625.520 800.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 796.000 652.400 800.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 796.000 679.280 800.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 796.000 706.160 800.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 796.000 733.040 800.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 796.000 759.920 800.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 796.000 786.800 800.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 796.000 813.680 800.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 796.000 840.560 800.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 796.000 114.800 800.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 796.000 867.440 800.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 893.760 796.000 894.320 800.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 920.640 796.000 921.200 800.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 796.000 948.080 800.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 796.000 974.960 800.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1001.280 796.000 1001.840 800.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 796.000 1028.720 800.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 796.000 1055.600 800.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 796.000 141.680 800.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 796.000 168.560 800.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 796.000 195.440 800.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 796.000 222.320 800.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 796.000 249.200 800.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 796.000 276.080 800.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 796.000 302.960 800.000 ;
    END
  END io_out[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 0.000 28.560 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 0.000 213.360 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 0.000 246.960 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 0.000 314.160 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 0.000 330.960 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 0.000 45.360 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 0.000 381.360 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 0.000 398.160 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 0.000 431.760 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 0.000 448.560 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 0.000 465.360 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 0.000 498.960 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 0.000 515.760 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 0.000 549.360 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 0.000 566.160 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 582.400 0.000 582.960 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 0.000 599.760 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 616.000 0.000 616.560 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 632.800 0.000 633.360 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 0.000 650.160 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 666.400 0.000 666.960 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 0.000 683.760 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 700.000 0.000 700.560 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 716.800 0.000 717.360 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 733.600 0.000 734.160 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 750.400 0.000 750.960 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 0.000 767.760 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 784.000 0.000 784.560 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 800.800 0.000 801.360 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 817.600 0.000 818.160 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 834.400 0.000 834.960 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 851.200 0.000 851.760 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 868.000 0.000 868.560 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 884.800 0.000 885.360 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 901.600 0.000 902.160 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 918.400 0.000 918.960 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 935.200 0.000 935.760 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 952.000 0.000 952.560 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 968.800 0.000 969.360 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 985.600 0.000 986.160 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1002.400 0.000 1002.960 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1019.200 0.000 1019.760 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1036.000 0.000 1036.560 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1052.800 0.000 1053.360 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1069.600 0.000 1070.160 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1086.400 0.000 1086.960 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END la_data_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 11.200 0.000 11.760 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 782.240 1093.550 784.430 ;
      LAYER Nwell ;
        RECT 6.290 777.920 1093.550 782.240 ;
      LAYER Pwell ;
        RECT 6.290 774.400 1093.550 777.920 ;
      LAYER Nwell ;
        RECT 6.290 770.080 1093.550 774.400 ;
      LAYER Pwell ;
        RECT 6.290 766.560 1093.550 770.080 ;
      LAYER Nwell ;
        RECT 6.290 762.240 1093.550 766.560 ;
      LAYER Pwell ;
        RECT 6.290 758.720 1093.550 762.240 ;
      LAYER Nwell ;
        RECT 6.290 754.400 1093.550 758.720 ;
      LAYER Pwell ;
        RECT 6.290 750.880 1093.550 754.400 ;
      LAYER Nwell ;
        RECT 6.290 746.560 1093.550 750.880 ;
      LAYER Pwell ;
        RECT 6.290 743.040 1093.550 746.560 ;
      LAYER Nwell ;
        RECT 6.290 738.720 1093.550 743.040 ;
      LAYER Pwell ;
        RECT 6.290 735.200 1093.550 738.720 ;
      LAYER Nwell ;
        RECT 6.290 730.880 1093.550 735.200 ;
      LAYER Pwell ;
        RECT 6.290 727.360 1093.550 730.880 ;
      LAYER Nwell ;
        RECT 6.290 727.235 292.360 727.360 ;
        RECT 6.290 723.165 1093.550 727.235 ;
        RECT 6.290 723.040 290.120 723.165 ;
      LAYER Pwell ;
        RECT 6.290 719.520 1093.550 723.040 ;
      LAYER Nwell ;
        RECT 6.290 719.395 266.600 719.520 ;
        RECT 6.290 715.325 1093.550 719.395 ;
        RECT 6.290 715.200 345.905 715.325 ;
      LAYER Pwell ;
        RECT 6.290 711.680 1093.550 715.200 ;
      LAYER Nwell ;
        RECT 6.290 711.555 260.785 711.680 ;
        RECT 6.290 707.485 1093.550 711.555 ;
        RECT 6.290 707.360 232.785 707.485 ;
      LAYER Pwell ;
        RECT 6.290 703.840 1093.550 707.360 ;
      LAYER Nwell ;
        RECT 6.290 703.715 227.745 703.840 ;
        RECT 6.290 699.645 1093.550 703.715 ;
        RECT 6.290 699.520 311.960 699.645 ;
      LAYER Pwell ;
        RECT 6.290 696.000 1093.550 699.520 ;
      LAYER Nwell ;
        RECT 6.290 695.875 210.385 696.000 ;
        RECT 6.290 691.805 1093.550 695.875 ;
        RECT 6.290 691.680 137.350 691.805 ;
      LAYER Pwell ;
        RECT 6.290 688.160 1093.550 691.680 ;
      LAYER Nwell ;
        RECT 6.290 688.035 188.310 688.160 ;
        RECT 6.290 683.965 1093.550 688.035 ;
        RECT 6.290 683.840 71.340 683.965 ;
      LAYER Pwell ;
        RECT 6.290 680.320 1093.550 683.840 ;
      LAYER Nwell ;
        RECT 6.290 680.195 69.460 680.320 ;
        RECT 6.290 676.125 1093.550 680.195 ;
        RECT 6.290 676.000 57.270 676.125 ;
      LAYER Pwell ;
        RECT 6.290 672.480 1093.550 676.000 ;
      LAYER Nwell ;
        RECT 6.290 672.355 175.430 672.480 ;
        RECT 6.290 668.285 1093.550 672.355 ;
        RECT 6.290 668.160 140.710 668.285 ;
      LAYER Pwell ;
        RECT 6.290 664.640 1093.550 668.160 ;
      LAYER Nwell ;
        RECT 6.290 664.515 57.270 664.640 ;
        RECT 6.290 660.445 1093.550 664.515 ;
        RECT 6.290 660.320 159.750 660.445 ;
      LAYER Pwell ;
        RECT 6.290 656.800 1093.550 660.320 ;
      LAYER Nwell ;
        RECT 6.290 656.675 185.230 656.800 ;
        RECT 6.290 652.605 1093.550 656.675 ;
        RECT 6.290 652.480 52.230 652.605 ;
      LAYER Pwell ;
        RECT 6.290 648.960 1093.550 652.480 ;
      LAYER Nwell ;
        RECT 6.290 648.835 36.865 648.960 ;
        RECT 6.290 644.765 1093.550 648.835 ;
        RECT 6.290 644.640 28.990 644.765 ;
      LAYER Pwell ;
        RECT 6.290 641.120 1093.550 644.640 ;
      LAYER Nwell ;
        RECT 6.290 640.995 117.470 641.120 ;
        RECT 6.290 636.925 1093.550 640.995 ;
        RECT 6.290 636.800 41.590 636.925 ;
      LAYER Pwell ;
        RECT 6.290 633.280 1093.550 636.800 ;
      LAYER Nwell ;
        RECT 6.290 633.155 34.870 633.280 ;
        RECT 6.290 629.085 1093.550 633.155 ;
        RECT 6.290 628.960 30.670 629.085 ;
      LAYER Pwell ;
        RECT 6.290 625.440 1093.550 628.960 ;
      LAYER Nwell ;
        RECT 6.290 625.315 66.510 625.440 ;
        RECT 6.290 621.245 1093.550 625.315 ;
        RECT 6.290 621.120 367.745 621.245 ;
      LAYER Pwell ;
        RECT 6.290 617.600 1093.550 621.120 ;
      LAYER Nwell ;
        RECT 6.290 617.475 160.870 617.600 ;
        RECT 6.290 613.405 1093.550 617.475 ;
        RECT 6.290 613.280 97.030 613.405 ;
      LAYER Pwell ;
        RECT 6.290 609.760 1093.550 613.280 ;
      LAYER Nwell ;
        RECT 6.290 609.635 156.715 609.760 ;
        RECT 6.290 605.565 1093.550 609.635 ;
        RECT 6.290 605.440 195.590 605.565 ;
      LAYER Pwell ;
        RECT 6.290 601.920 1093.550 605.440 ;
      LAYER Nwell ;
        RECT 6.290 601.795 301.195 601.920 ;
        RECT 6.290 597.725 1093.550 601.795 ;
        RECT 6.290 597.600 111.445 597.725 ;
      LAYER Pwell ;
        RECT 6.290 594.080 1093.550 597.600 ;
      LAYER Nwell ;
        RECT 6.290 593.955 110.470 594.080 ;
        RECT 6.290 589.885 1093.550 593.955 ;
        RECT 6.290 589.760 357.865 589.885 ;
      LAYER Pwell ;
        RECT 6.290 586.240 1093.550 589.760 ;
      LAYER Nwell ;
        RECT 6.290 586.115 236.540 586.240 ;
        RECT 6.290 582.045 1093.550 586.115 ;
        RECT 6.290 581.920 71.505 582.045 ;
      LAYER Pwell ;
        RECT 6.290 578.400 1093.550 581.920 ;
      LAYER Nwell ;
        RECT 6.290 578.275 101.960 578.400 ;
        RECT 6.290 574.205 1093.550 578.275 ;
        RECT 6.290 574.080 90.200 574.205 ;
      LAYER Pwell ;
        RECT 6.290 570.560 1093.550 574.080 ;
      LAYER Nwell ;
        RECT 6.290 570.435 58.840 570.560 ;
        RECT 6.290 566.365 1093.550 570.435 ;
        RECT 6.290 566.240 110.785 566.365 ;
      LAYER Pwell ;
        RECT 6.290 562.720 1093.550 566.240 ;
      LAYER Nwell ;
        RECT 6.290 562.595 92.785 562.720 ;
        RECT 6.290 558.525 1093.550 562.595 ;
        RECT 6.290 558.400 85.585 558.525 ;
      LAYER Pwell ;
        RECT 6.290 554.880 1093.550 558.400 ;
      LAYER Nwell ;
        RECT 6.290 554.755 59.745 554.880 ;
        RECT 6.290 550.685 1093.550 554.755 ;
        RECT 6.290 550.560 239.900 550.685 ;
      LAYER Pwell ;
        RECT 6.290 547.040 1093.550 550.560 ;
      LAYER Nwell ;
        RECT 6.290 546.915 129.275 547.040 ;
        RECT 6.290 542.845 1093.550 546.915 ;
        RECT 6.290 542.720 110.120 542.845 ;
      LAYER Pwell ;
        RECT 6.290 539.200 1093.550 542.720 ;
      LAYER Nwell ;
        RECT 6.290 539.075 147.245 539.200 ;
        RECT 6.290 535.005 1093.550 539.075 ;
        RECT 6.290 534.880 51.905 535.005 ;
      LAYER Pwell ;
        RECT 6.290 531.360 1093.550 534.880 ;
      LAYER Nwell ;
        RECT 6.290 531.235 139.450 531.360 ;
        RECT 6.290 527.165 1093.550 531.235 ;
        RECT 6.290 527.040 46.520 527.165 ;
      LAYER Pwell ;
        RECT 6.290 523.520 1093.550 527.040 ;
      LAYER Nwell ;
        RECT 6.290 523.395 71.550 523.520 ;
        RECT 6.290 519.325 1093.550 523.395 ;
        RECT 6.290 519.200 122.555 519.325 ;
      LAYER Pwell ;
        RECT 6.290 515.680 1093.550 519.200 ;
      LAYER Nwell ;
        RECT 6.290 515.555 72.825 515.680 ;
        RECT 6.290 511.485 1093.550 515.555 ;
        RECT 6.290 511.360 174.380 511.485 ;
      LAYER Pwell ;
        RECT 6.290 507.840 1093.550 511.360 ;
      LAYER Nwell ;
        RECT 6.290 507.715 66.035 507.840 ;
        RECT 6.290 503.645 1093.550 507.715 ;
        RECT 6.290 503.520 60.385 503.645 ;
      LAYER Pwell ;
        RECT 6.290 500.000 1093.550 503.520 ;
      LAYER Nwell ;
        RECT 6.290 499.875 96.225 500.000 ;
        RECT 6.290 495.805 1093.550 499.875 ;
        RECT 6.290 495.680 67.780 495.805 ;
      LAYER Pwell ;
        RECT 6.290 492.160 1093.550 495.680 ;
      LAYER Nwell ;
        RECT 6.290 492.035 153.915 492.160 ;
        RECT 6.290 487.965 1093.550 492.035 ;
        RECT 6.290 487.840 56.450 487.965 ;
      LAYER Pwell ;
        RECT 6.290 484.320 1093.550 487.840 ;
      LAYER Nwell ;
        RECT 6.290 484.195 96.185 484.320 ;
        RECT 6.290 480.125 1093.550 484.195 ;
        RECT 6.290 480.000 475.980 480.125 ;
      LAYER Pwell ;
        RECT 6.290 476.480 1093.550 480.000 ;
      LAYER Nwell ;
        RECT 6.290 476.355 76.310 476.480 ;
        RECT 6.290 472.285 1093.550 476.355 ;
        RECT 6.290 472.160 501.115 472.285 ;
      LAYER Pwell ;
        RECT 6.290 468.640 1093.550 472.160 ;
      LAYER Nwell ;
        RECT 6.290 468.515 102.070 468.640 ;
        RECT 6.290 464.445 1093.550 468.515 ;
        RECT 6.290 464.320 190.355 464.445 ;
      LAYER Pwell ;
        RECT 6.290 460.800 1093.550 464.320 ;
      LAYER Nwell ;
        RECT 6.290 460.675 101.745 460.800 ;
        RECT 6.290 456.605 1093.550 460.675 ;
        RECT 6.290 456.480 522.995 456.605 ;
      LAYER Pwell ;
        RECT 6.290 452.960 1093.550 456.480 ;
      LAYER Nwell ;
        RECT 6.290 452.835 63.105 452.960 ;
        RECT 6.290 448.765 1093.550 452.835 ;
        RECT 6.290 448.640 168.650 448.765 ;
      LAYER Pwell ;
        RECT 6.290 445.120 1093.550 448.640 ;
      LAYER Nwell ;
        RECT 6.290 444.995 70.040 445.120 ;
        RECT 6.290 440.925 1093.550 444.995 ;
        RECT 6.290 440.800 237.980 440.925 ;
      LAYER Pwell ;
        RECT 6.290 437.280 1093.550 440.800 ;
      LAYER Nwell ;
        RECT 6.290 437.155 98.385 437.280 ;
        RECT 6.290 433.085 1093.550 437.155 ;
        RECT 6.290 432.960 71.505 433.085 ;
      LAYER Pwell ;
        RECT 6.290 429.440 1093.550 432.960 ;
      LAYER Nwell ;
        RECT 6.290 429.315 61.985 429.440 ;
        RECT 6.290 425.245 1093.550 429.315 ;
        RECT 6.290 425.120 187.555 425.245 ;
      LAYER Pwell ;
        RECT 6.290 421.600 1093.550 425.120 ;
      LAYER Nwell ;
        RECT 6.290 421.475 187.465 421.600 ;
        RECT 6.290 417.405 1093.550 421.475 ;
        RECT 6.290 417.280 81.585 417.405 ;
      LAYER Pwell ;
        RECT 6.290 413.760 1093.550 417.280 ;
      LAYER Nwell ;
        RECT 6.290 413.635 185.785 413.760 ;
        RECT 6.290 409.565 1093.550 413.635 ;
        RECT 6.290 409.440 131.640 409.565 ;
      LAYER Pwell ;
        RECT 6.290 405.920 1093.550 409.440 ;
      LAYER Nwell ;
        RECT 6.290 405.795 103.640 405.920 ;
        RECT 6.290 401.725 1093.550 405.795 ;
        RECT 6.290 401.600 110.705 401.725 ;
      LAYER Pwell ;
        RECT 6.290 398.080 1093.550 401.600 ;
      LAYER Nwell ;
        RECT 6.290 397.955 183.605 398.080 ;
        RECT 6.290 393.885 1093.550 397.955 ;
        RECT 6.290 393.760 132.200 393.885 ;
      LAYER Pwell ;
        RECT 6.290 390.240 1093.550 393.760 ;
      LAYER Nwell ;
        RECT 6.290 390.115 366.105 390.240 ;
        RECT 6.290 386.045 1093.550 390.115 ;
        RECT 6.290 385.920 123.240 386.045 ;
      LAYER Pwell ;
        RECT 6.290 382.400 1093.550 385.920 ;
      LAYER Nwell ;
        RECT 6.290 382.275 142.625 382.400 ;
        RECT 6.290 378.205 1093.550 382.275 ;
        RECT 6.290 378.080 128.625 378.205 ;
      LAYER Pwell ;
        RECT 6.290 374.560 1093.550 378.080 ;
      LAYER Nwell ;
        RECT 6.290 374.435 256.865 374.560 ;
        RECT 6.290 370.365 1093.550 374.435 ;
        RECT 6.290 370.240 123.585 370.365 ;
      LAYER Pwell ;
        RECT 6.290 366.720 1093.550 370.240 ;
      LAYER Nwell ;
        RECT 6.290 366.595 186.865 366.720 ;
        RECT 6.290 362.525 1093.550 366.595 ;
        RECT 6.290 362.400 136.120 362.525 ;
      LAYER Pwell ;
        RECT 6.290 358.880 1093.550 362.400 ;
      LAYER Nwell ;
        RECT 6.290 358.755 148.785 358.880 ;
        RECT 6.290 354.685 1093.550 358.755 ;
        RECT 6.290 354.560 120.225 354.685 ;
      LAYER Pwell ;
        RECT 6.290 351.040 1093.550 354.560 ;
      LAYER Nwell ;
        RECT 6.290 350.915 141.720 351.040 ;
        RECT 6.290 346.845 1093.550 350.915 ;
        RECT 6.290 346.720 95.800 346.845 ;
      LAYER Pwell ;
        RECT 6.290 343.200 1093.550 346.720 ;
      LAYER Nwell ;
        RECT 6.290 343.075 111.825 343.200 ;
        RECT 6.290 339.005 1093.550 343.075 ;
        RECT 6.290 338.880 71.505 339.005 ;
      LAYER Pwell ;
        RECT 6.290 335.360 1093.550 338.880 ;
      LAYER Nwell ;
        RECT 6.290 335.235 61.425 335.360 ;
        RECT 6.290 331.165 1093.550 335.235 ;
        RECT 6.290 331.040 61.555 331.165 ;
      LAYER Pwell ;
        RECT 6.290 327.520 1093.550 331.040 ;
      LAYER Nwell ;
        RECT 6.290 327.395 55.395 327.520 ;
        RECT 6.290 323.325 1093.550 327.395 ;
        RECT 6.290 323.200 49.320 323.325 ;
      LAYER Pwell ;
        RECT 6.290 319.680 1093.550 323.200 ;
      LAYER Nwell ;
        RECT 6.290 319.555 91.105 319.680 ;
        RECT 6.290 315.485 1093.550 319.555 ;
        RECT 6.290 315.360 42.385 315.485 ;
      LAYER Pwell ;
        RECT 6.290 311.840 1093.550 315.360 ;
      LAYER Nwell ;
        RECT 6.290 307.645 1093.550 311.840 ;
        RECT 6.290 307.520 198.630 307.645 ;
      LAYER Pwell ;
        RECT 6.290 304.000 1093.550 307.520 ;
      LAYER Nwell ;
        RECT 6.290 303.875 63.665 304.000 ;
        RECT 6.290 299.805 1093.550 303.875 ;
        RECT 6.290 299.680 123.025 299.805 ;
      LAYER Pwell ;
        RECT 6.290 296.160 1093.550 299.680 ;
      LAYER Nwell ;
        RECT 6.290 296.035 21.105 296.160 ;
        RECT 6.290 291.965 1093.550 296.035 ;
        RECT 6.290 291.840 13.825 291.965 ;
      LAYER Pwell ;
        RECT 6.290 288.320 1093.550 291.840 ;
      LAYER Nwell ;
        RECT 6.290 288.195 14.945 288.320 ;
        RECT 6.290 284.125 1093.550 288.195 ;
        RECT 6.290 284.000 84.385 284.125 ;
      LAYER Pwell ;
        RECT 6.290 280.480 1093.550 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 423.400 280.480 ;
        RECT 6.290 276.285 1093.550 280.355 ;
        RECT 6.290 276.160 78.785 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 1093.550 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 18.305 272.640 ;
        RECT 6.290 268.445 1093.550 272.515 ;
        RECT 6.290 268.320 32.305 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 1093.550 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 150.465 264.800 ;
        RECT 6.290 260.605 1093.550 264.675 ;
        RECT 6.290 260.480 14.945 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 1093.550 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 20.545 256.960 ;
        RECT 6.290 252.765 1093.550 256.835 ;
        RECT 6.290 252.640 78.785 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 1093.550 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 18.305 249.120 ;
        RECT 6.290 244.925 1093.550 248.995 ;
        RECT 6.290 244.800 14.945 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 1093.550 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 353.400 241.280 ;
        RECT 6.290 237.085 1093.550 241.155 ;
        RECT 6.290 236.960 76.545 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 1093.550 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 149.345 233.440 ;
        RECT 6.290 229.245 1093.550 233.315 ;
        RECT 6.290 229.120 13.825 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 1093.550 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 18.865 225.600 ;
        RECT 6.290 221.405 1093.550 225.475 ;
        RECT 6.290 221.280 54.920 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 1093.550 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 25.585 217.760 ;
        RECT 6.290 213.565 1093.550 217.635 ;
        RECT 6.290 213.440 85.505 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 1093.550 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 151.025 209.920 ;
        RECT 6.290 205.725 1093.550 209.795 ;
        RECT 6.290 205.600 123.585 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 1093.550 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 20.545 202.080 ;
        RECT 6.290 197.885 1093.550 201.955 ;
        RECT 6.290 197.760 189.105 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 1093.550 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 217.320 194.240 ;
        RECT 6.290 190.045 1093.550 194.115 ;
        RECT 6.290 189.920 14.945 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 1093.550 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 53.585 186.400 ;
        RECT 6.290 182.205 1093.550 186.275 ;
        RECT 6.290 182.080 158.305 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 1093.550 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 19.985 178.560 ;
        RECT 6.290 174.365 1093.550 178.435 ;
        RECT 6.290 174.240 238.035 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 1093.550 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 21.105 170.720 ;
        RECT 6.290 166.525 1093.550 170.595 ;
        RECT 6.290 166.400 32.305 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 1093.550 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 26.920 162.880 ;
        RECT 6.290 158.685 1093.550 162.755 ;
        RECT 6.290 158.560 231.105 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 1093.550 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 190.225 155.040 ;
        RECT 6.290 150.845 1093.550 154.915 ;
        RECT 6.290 150.720 37.345 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 1093.550 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 59.185 147.200 ;
        RECT 6.290 143.005 1093.550 147.075 ;
        RECT 6.290 142.880 54.145 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 1093.550 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 54.145 139.360 ;
        RECT 6.290 135.165 1093.550 139.235 ;
        RECT 6.290 135.040 215.080 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 1093.550 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 118.200 131.520 ;
        RECT 6.290 127.325 1093.550 131.395 ;
        RECT 6.290 127.200 156.065 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 1093.550 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 223.825 123.680 ;
        RECT 6.290 119.485 1093.550 123.555 ;
        RECT 6.290 119.360 129.745 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 1093.550 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 339.400 115.840 ;
        RECT 6.290 111.645 1093.550 115.715 ;
        RECT 6.290 111.520 132.545 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 1093.550 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 292.705 108.000 ;
        RECT 6.290 103.805 1093.550 107.875 ;
        RECT 6.290 103.680 163.905 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 1093.550 103.680 ;
      LAYER Nwell ;
        RECT 6.290 95.965 1093.550 100.160 ;
        RECT 6.290 95.840 163.905 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 1093.550 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 216.545 92.320 ;
        RECT 6.290 88.125 1093.550 92.195 ;
        RECT 6.290 88.000 236.705 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 1093.550 88.000 ;
      LAYER Nwell ;
        RECT 6.290 80.160 1093.550 84.480 ;
      LAYER Pwell ;
        RECT 6.290 76.640 1093.550 80.160 ;
      LAYER Nwell ;
        RECT 6.290 72.320 1093.550 76.640 ;
      LAYER Pwell ;
        RECT 6.290 68.800 1093.550 72.320 ;
      LAYER Nwell ;
        RECT 6.290 64.480 1093.550 68.800 ;
      LAYER Pwell ;
        RECT 6.290 60.960 1093.550 64.480 ;
      LAYER Nwell ;
        RECT 6.290 56.640 1093.550 60.960 ;
      LAYER Pwell ;
        RECT 6.290 53.120 1093.550 56.640 ;
      LAYER Nwell ;
        RECT 6.290 48.800 1093.550 53.120 ;
      LAYER Pwell ;
        RECT 6.290 45.280 1093.550 48.800 ;
      LAYER Nwell ;
        RECT 6.290 40.960 1093.550 45.280 ;
      LAYER Pwell ;
        RECT 6.290 37.440 1093.550 40.960 ;
      LAYER Nwell ;
        RECT 6.290 33.120 1093.550 37.440 ;
      LAYER Pwell ;
        RECT 6.290 29.600 1093.550 33.120 ;
      LAYER Nwell ;
        RECT 6.290 25.280 1093.550 29.600 ;
      LAYER Pwell ;
        RECT 6.290 21.760 1093.550 25.280 ;
      LAYER Nwell ;
        RECT 6.290 17.440 1093.550 21.760 ;
      LAYER Pwell ;
        RECT 6.290 15.250 1093.550 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1093.120 786.090 ;
      LAYER Metal2 ;
        RECT 7.980 795.700 42.260 796.740 ;
        RECT 43.420 795.700 51.220 796.740 ;
        RECT 52.380 795.700 60.180 796.740 ;
        RECT 61.340 795.700 69.140 796.740 ;
        RECT 70.300 795.700 78.100 796.740 ;
        RECT 79.260 795.700 87.060 796.740 ;
        RECT 88.220 795.700 96.020 796.740 ;
        RECT 97.180 795.700 104.980 796.740 ;
        RECT 106.140 795.700 113.940 796.740 ;
        RECT 115.100 795.700 122.900 796.740 ;
        RECT 124.060 795.700 131.860 796.740 ;
        RECT 133.020 795.700 140.820 796.740 ;
        RECT 141.980 795.700 149.780 796.740 ;
        RECT 150.940 795.700 158.740 796.740 ;
        RECT 159.900 795.700 167.700 796.740 ;
        RECT 168.860 795.700 176.660 796.740 ;
        RECT 177.820 795.700 185.620 796.740 ;
        RECT 186.780 795.700 194.580 796.740 ;
        RECT 195.740 795.700 203.540 796.740 ;
        RECT 204.700 795.700 212.500 796.740 ;
        RECT 213.660 795.700 221.460 796.740 ;
        RECT 222.620 795.700 230.420 796.740 ;
        RECT 231.580 795.700 239.380 796.740 ;
        RECT 240.540 795.700 248.340 796.740 ;
        RECT 249.500 795.700 257.300 796.740 ;
        RECT 258.460 795.700 266.260 796.740 ;
        RECT 267.420 795.700 275.220 796.740 ;
        RECT 276.380 795.700 284.180 796.740 ;
        RECT 285.340 795.700 293.140 796.740 ;
        RECT 294.300 795.700 302.100 796.740 ;
        RECT 303.260 795.700 311.060 796.740 ;
        RECT 312.220 795.700 320.020 796.740 ;
        RECT 321.180 795.700 328.980 796.740 ;
        RECT 330.140 795.700 337.940 796.740 ;
        RECT 339.100 795.700 346.900 796.740 ;
        RECT 348.060 795.700 355.860 796.740 ;
        RECT 357.020 795.700 364.820 796.740 ;
        RECT 365.980 795.700 373.780 796.740 ;
        RECT 374.940 795.700 382.740 796.740 ;
        RECT 383.900 795.700 391.700 796.740 ;
        RECT 392.860 795.700 400.660 796.740 ;
        RECT 401.820 795.700 409.620 796.740 ;
        RECT 410.780 795.700 418.580 796.740 ;
        RECT 419.740 795.700 427.540 796.740 ;
        RECT 428.700 795.700 436.500 796.740 ;
        RECT 437.660 795.700 445.460 796.740 ;
        RECT 446.620 795.700 454.420 796.740 ;
        RECT 455.580 795.700 463.380 796.740 ;
        RECT 464.540 795.700 472.340 796.740 ;
        RECT 473.500 795.700 481.300 796.740 ;
        RECT 482.460 795.700 490.260 796.740 ;
        RECT 491.420 795.700 499.220 796.740 ;
        RECT 500.380 795.700 508.180 796.740 ;
        RECT 509.340 795.700 517.140 796.740 ;
        RECT 518.300 795.700 526.100 796.740 ;
        RECT 527.260 795.700 535.060 796.740 ;
        RECT 536.220 795.700 544.020 796.740 ;
        RECT 545.180 795.700 552.980 796.740 ;
        RECT 554.140 795.700 561.940 796.740 ;
        RECT 563.100 795.700 570.900 796.740 ;
        RECT 572.060 795.700 579.860 796.740 ;
        RECT 581.020 795.700 588.820 796.740 ;
        RECT 589.980 795.700 597.780 796.740 ;
        RECT 598.940 795.700 606.740 796.740 ;
        RECT 607.900 795.700 615.700 796.740 ;
        RECT 616.860 795.700 624.660 796.740 ;
        RECT 625.820 795.700 633.620 796.740 ;
        RECT 634.780 795.700 642.580 796.740 ;
        RECT 643.740 795.700 651.540 796.740 ;
        RECT 652.700 795.700 660.500 796.740 ;
        RECT 661.660 795.700 669.460 796.740 ;
        RECT 670.620 795.700 678.420 796.740 ;
        RECT 679.580 795.700 687.380 796.740 ;
        RECT 688.540 795.700 696.340 796.740 ;
        RECT 697.500 795.700 705.300 796.740 ;
        RECT 706.460 795.700 714.260 796.740 ;
        RECT 715.420 795.700 723.220 796.740 ;
        RECT 724.380 795.700 732.180 796.740 ;
        RECT 733.340 795.700 741.140 796.740 ;
        RECT 742.300 795.700 750.100 796.740 ;
        RECT 751.260 795.700 759.060 796.740 ;
        RECT 760.220 795.700 768.020 796.740 ;
        RECT 769.180 795.700 776.980 796.740 ;
        RECT 778.140 795.700 785.940 796.740 ;
        RECT 787.100 795.700 794.900 796.740 ;
        RECT 796.060 795.700 803.860 796.740 ;
        RECT 805.020 795.700 812.820 796.740 ;
        RECT 813.980 795.700 821.780 796.740 ;
        RECT 822.940 795.700 830.740 796.740 ;
        RECT 831.900 795.700 839.700 796.740 ;
        RECT 840.860 795.700 848.660 796.740 ;
        RECT 849.820 795.700 857.620 796.740 ;
        RECT 858.780 795.700 866.580 796.740 ;
        RECT 867.740 795.700 875.540 796.740 ;
        RECT 876.700 795.700 884.500 796.740 ;
        RECT 885.660 795.700 893.460 796.740 ;
        RECT 894.620 795.700 902.420 796.740 ;
        RECT 903.580 795.700 911.380 796.740 ;
        RECT 912.540 795.700 920.340 796.740 ;
        RECT 921.500 795.700 929.300 796.740 ;
        RECT 930.460 795.700 938.260 796.740 ;
        RECT 939.420 795.700 947.220 796.740 ;
        RECT 948.380 795.700 956.180 796.740 ;
        RECT 957.340 795.700 965.140 796.740 ;
        RECT 966.300 795.700 974.100 796.740 ;
        RECT 975.260 795.700 983.060 796.740 ;
        RECT 984.220 795.700 992.020 796.740 ;
        RECT 993.180 795.700 1000.980 796.740 ;
        RECT 1002.140 795.700 1009.940 796.740 ;
        RECT 1011.100 795.700 1018.900 796.740 ;
        RECT 1020.060 795.700 1027.860 796.740 ;
        RECT 1029.020 795.700 1036.820 796.740 ;
        RECT 1037.980 795.700 1045.780 796.740 ;
        RECT 1046.940 795.700 1054.740 796.740 ;
        RECT 1055.900 795.700 1087.940 796.740 ;
        RECT 7.980 4.300 1087.940 795.700 ;
        RECT 7.980 3.500 10.900 4.300 ;
        RECT 12.060 3.500 27.700 4.300 ;
        RECT 28.860 3.500 44.500 4.300 ;
        RECT 45.660 3.500 61.300 4.300 ;
        RECT 62.460 3.500 78.100 4.300 ;
        RECT 79.260 3.500 94.900 4.300 ;
        RECT 96.060 3.500 111.700 4.300 ;
        RECT 112.860 3.500 128.500 4.300 ;
        RECT 129.660 3.500 145.300 4.300 ;
        RECT 146.460 3.500 162.100 4.300 ;
        RECT 163.260 3.500 178.900 4.300 ;
        RECT 180.060 3.500 195.700 4.300 ;
        RECT 196.860 3.500 212.500 4.300 ;
        RECT 213.660 3.500 229.300 4.300 ;
        RECT 230.460 3.500 246.100 4.300 ;
        RECT 247.260 3.500 262.900 4.300 ;
        RECT 264.060 3.500 279.700 4.300 ;
        RECT 280.860 3.500 296.500 4.300 ;
        RECT 297.660 3.500 313.300 4.300 ;
        RECT 314.460 3.500 330.100 4.300 ;
        RECT 331.260 3.500 346.900 4.300 ;
        RECT 348.060 3.500 363.700 4.300 ;
        RECT 364.860 3.500 380.500 4.300 ;
        RECT 381.660 3.500 397.300 4.300 ;
        RECT 398.460 3.500 414.100 4.300 ;
        RECT 415.260 3.500 430.900 4.300 ;
        RECT 432.060 3.500 447.700 4.300 ;
        RECT 448.860 3.500 464.500 4.300 ;
        RECT 465.660 3.500 481.300 4.300 ;
        RECT 482.460 3.500 498.100 4.300 ;
        RECT 499.260 3.500 514.900 4.300 ;
        RECT 516.060 3.500 531.700 4.300 ;
        RECT 532.860 3.500 548.500 4.300 ;
        RECT 549.660 3.500 565.300 4.300 ;
        RECT 566.460 3.500 582.100 4.300 ;
        RECT 583.260 3.500 598.900 4.300 ;
        RECT 600.060 3.500 615.700 4.300 ;
        RECT 616.860 3.500 632.500 4.300 ;
        RECT 633.660 3.500 649.300 4.300 ;
        RECT 650.460 3.500 666.100 4.300 ;
        RECT 667.260 3.500 682.900 4.300 ;
        RECT 684.060 3.500 699.700 4.300 ;
        RECT 700.860 3.500 716.500 4.300 ;
        RECT 717.660 3.500 733.300 4.300 ;
        RECT 734.460 3.500 750.100 4.300 ;
        RECT 751.260 3.500 766.900 4.300 ;
        RECT 768.060 3.500 783.700 4.300 ;
        RECT 784.860 3.500 800.500 4.300 ;
        RECT 801.660 3.500 817.300 4.300 ;
        RECT 818.460 3.500 834.100 4.300 ;
        RECT 835.260 3.500 850.900 4.300 ;
        RECT 852.060 3.500 867.700 4.300 ;
        RECT 868.860 3.500 884.500 4.300 ;
        RECT 885.660 3.500 901.300 4.300 ;
        RECT 902.460 3.500 918.100 4.300 ;
        RECT 919.260 3.500 934.900 4.300 ;
        RECT 936.060 3.500 951.700 4.300 ;
        RECT 952.860 3.500 968.500 4.300 ;
        RECT 969.660 3.500 985.300 4.300 ;
        RECT 986.460 3.500 1002.100 4.300 ;
        RECT 1003.260 3.500 1018.900 4.300 ;
        RECT 1020.060 3.500 1035.700 4.300 ;
        RECT 1036.860 3.500 1052.500 4.300 ;
        RECT 1053.660 3.500 1069.300 4.300 ;
        RECT 1070.460 3.500 1086.100 4.300 ;
        RECT 1087.260 3.500 1087.940 4.300 ;
      LAYER Metal3 ;
        RECT 7.930 5.180 1022.150 793.380 ;
      LAYER Metal4 ;
        RECT 51.100 784.600 773.220 793.430 ;
        RECT 51.100 15.080 98.740 784.600 ;
        RECT 100.940 15.080 175.540 784.600 ;
        RECT 177.740 15.080 252.340 784.600 ;
        RECT 254.540 15.080 329.140 784.600 ;
        RECT 331.340 15.080 405.940 784.600 ;
        RECT 408.140 15.080 482.740 784.600 ;
        RECT 484.940 15.080 559.540 784.600 ;
        RECT 561.740 15.080 636.340 784.600 ;
        RECT 638.540 15.080 713.140 784.600 ;
        RECT 715.340 15.080 773.220 784.600 ;
        RECT 51.100 5.130 773.220 15.080 ;
  END
END wrapped_as2650
END LIBRARY

