* NGSPICE file created from serial_ports.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

.subckt serial_ports RXD TXD addr[0] addr[1] addr[2] bus_cyc bus_we data_in[0] data_in[1]
+ data_in[2] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7] data_out[0] data_out[1]
+ data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] io_in io_oeb[0]
+ io_oeb[1] io_oeb[2] io_out[0] io_out[1] irq3 rst vdd vss wb_clk_i io_out[2]
XFILLER_0_49_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1206__A1 _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1724__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1270_ _0615_ _0616_ uart.receiving _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1606_ _0432_ _0568_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0985_ spi.div_counter\[4\] _0379_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1537_ _0816_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1399_ uart.div_counter\[2\] uart.divisor\[2\] _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1468_ _0780_ _0781_ _0783_ _0574_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1747__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1418__A1 uart.div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1322_ _0659_ _0661_ _0629_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1253_ _0253_ _0599_ _0604_ _0430_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1184_ _0527_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0968_ _0367_ _0361_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0899_ spi.data_out_buff\[3\] _0306_ _0311_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_2_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0871__A2 spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0836__I spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1305_ _0617_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1236_ uart.divisor\[15\] _0576_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1167_ uart.receive_div_counter\[11\] uart.divisor\[11\] _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1098_ _0286_ _0275_ _0473_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_19_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1021_ _0408_ _0409_ _0411_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1785_ _0125_ clknet_4_11_0_wb_clk_i uart.has_byte vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1219_ uart.divisor\[10\] _0577_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_27_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1570_ _0179_ _0181_ _0169_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1780__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1004_ _0397_ _0398_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1768_ _0108_ clknet_4_1_0_wb_clk_i uart.data_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1699_ _0039_ clknet_4_9_0_wb_clk_i uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_12_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 data_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1527__A3 uart.div_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1622_ spi.data_in_buff\[3\] _0218_ _0221_ spi.data_in_buff\[4\] _0222_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1553_ uart.div_counter\[7\] _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1484_ _0793_ _0781_ _0796_ _0792_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_49_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1454__A2 _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1676__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1390__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1142__A1 uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0956__A1 spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1699__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0984_ spi.div_counter\[5\] _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1605_ _0209_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1536_ uart.div_counter\[4\] _0152_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1398_ _0719_ uart.divisor\[15\] _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1467_ uart.data_buff\[1\] _0768_ _0777_ _0782_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_60_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1418__A2 uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1321_ _0660_ _0626_ _0654_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1252_ _0440_ _0603_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1183_ uart.receive_counter\[0\] _0550_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1349__B _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0967_ _0368_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1714__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1519_ _0820_ _0824_ _0779_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0898_ _0308_ _0309_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0942__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1737__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1304_ uart.receive_div_counter\[4\] _0646_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1166_ uart.receive_div_counter\[1\] uart.divisor\[1\] _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1235_ _0454_ _0584_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1097_ net2 _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1020_ _0410_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1784_ _0124_ clknet_4_4_0_wb_clk_i uart.div_counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1218_ _0437_ _0571_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1149_ uart.divisor\[6\] _0507_ _0479_ spi.divisor\[6\] _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_27_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1003__A3 _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1003_ _0335_ spi.data_out_buff\[7\] _0349_ _0337_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_16_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1698_ _0038_ clknet_4_9_0_wb_clk_i uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1767_ _0107_ clknet_4_1_0_wb_clk_i uart.data_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input11_I data_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput21 net21 data_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1527__A4 uart.div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1160__A2 uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1552_ uart.div_counter\[7\] _0162_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1621_ _0214_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input3_I addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1483_ _0440_ _0794_ _0789_ _0795_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_43_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1770__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0956__A2 _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1016__I _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0947__A2 _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0983_ _0318_ _0381_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1604_ _0716_ _0699_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1635__B _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1535_ _0148_ _0150_ _0151_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1397_ uart.div_counter\[15\] _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1466_ _0280_ _0746_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1060__A1 uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1793__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1320_ uart.receive_div_counter\[7\] _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1051__A1 _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1182_ _0527_ _0538_ _0549_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1251_ _0598_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1666__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1042__A1 _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0897_ _0271_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0966_ _0314_ _0351_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1518_ _0821_ _0812_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_2_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1449_ _0746_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1303_ _0618_ _0644_ _0645_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_24_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1165_ uart.receive_div_counter\[13\] uart.divisor\[13\] _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1096_ _0460_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1234_ _0589_ _0590_ _0583_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0838__B2 spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0838__A1 spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1263__A1 spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0949_ _0344_ _0352_ _0340_ spi.counter\[4\] _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_38_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1254__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1006__A1 spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1493__A1 _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1783_ _0123_ clknet_4_4_0_wb_clk_i uart.div_counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1217_ _0575_ _0578_ _0420_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1079_ _0447_ _0455_ _0456_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1148_ spi.dout\[6\] _0499_ _0505_ uart.divisor\[14\] _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_27_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1236__A1 uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1727__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1019__I _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1463__B _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1002_ _0296_ _0376_ _0396_ net27 _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1466__A1 _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1218__A1 _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1697_ _0037_ clknet_4_9_0_wb_clk_i uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1766_ _0106_ clknet_4_1_0_wb_clk_i uart.data_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1209__A1 uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput22 net22 data_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1551_ _0163_ _0165_ _0779_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1620_ _0216_ _0220_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1482_ _0788_ _0785_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1749_ _0089_ clknet_4_15_0_wb_clk_i uart.receive_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1127__B1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1188__B _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0982_ spi.div_counter\[4\] _0369_ _0376_ _0380_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1109__B1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1603_ _0204_ _0207_ _0208_ _0719_ _0765_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1534_ _0746_ _0752_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1465_ _0774_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1396_ _0642_ _0614_ _0718_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0883__A2 _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1181_ _0543_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1250_ _0258_ _0599_ _0602_ _0430_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0896_ net11 _0290_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0965_ spi.div_counter\[1\] _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1517_ _0822_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1448_ _0764_ _0766_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1379_ uart.receive_buff\[2\] _0702_ _0704_ uart.receive_buff\[3\] _0708_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_2_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1760__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1302_ _0552_ net1 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1233_ uart.divisor\[14\] _0576_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1164_ _0528_ _0529_ _0530_ _0531_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1095_ _0466_ _0470_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1783__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0948_ _0344_ spi.counter\[4\] _0352_ _0340_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0879_ _0285_ _0294_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1305__I _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1040__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1782_ _0122_ clknet_4_5_0_wb_clk_i uart.div_counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1216_ uart.divisor\[9\] _0577_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1147_ uart.dout\[6\] _0465_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1078_ uart.divisor\[7\] _0445_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1679__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0874__I _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1001_ _0395_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1466__A2 _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1765_ _0105_ clknet_4_3_0_wb_clk_i uart.data_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1696_ _0036_ clknet_4_12_0_wb_clk_i uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__1154__B2 uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput23 net23 data_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1550_ _0156_ _0150_ _0164_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_34_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1136__A1 uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1481_ _0759_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1136__B2 spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1748_ _0088_ clknet_4_15_0_wb_clk_i uart.receive_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1127__A1 spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1679_ _0019_ clknet_4_2_0_wb_clk_i spi.div_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0981_ spi.div_counter\[4\] _0379_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1602_ uart.div_counter\[14\] _0827_ _0205_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1395_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1109__A1 uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1109__B2 uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1533_ _0149_ _0146_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1464_ uart.data_buff\[2\] _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1133__I _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1308__I _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1180_ _0544_ _0545_ _0546_ _0547_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__0882__I _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0964_ _0361_ _0362_ _0365_ _0366_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_54_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1516_ _0754_ _0752_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0895_ spi.data_out_buff\[4\] _0307_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1378_ _0458_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1502__A1 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1447_ uart.counter\[2\] _0749_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1038__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1301_ _0643_ _0640_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1232_ _0451_ _0584_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1163_ uart.receive_div_counter\[10\] uart.divisor\[10\] _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1094_ uart_ien _0467_ _0469_ uart.divisor\[8\] _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0947_ _0350_ _0351_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0878_ spi.data_out_buff\[0\] _0272_ _0293_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_13_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1781_ _0121_ clknet_4_5_0_wb_clk_i uart.div_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1750__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1146_ _0458_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1215_ _0576_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1077_ _0454_ _0433_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1172__A2 uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1773__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1163__A2 uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1000_ _0394_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1764_ _0104_ clknet_4_0_0_wb_clk_i uart.data_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1695_ _0035_ clknet_4_12_0_wb_clk_i uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1129_ _0472_ _0498_ _0500_ _0501_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1796__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1090__A1 uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 data_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1393__A2 _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0959__A2 _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1480_ uart.data_buff\[5\] _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1669__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1747_ _0087_ clknet_4_13_0_wb_clk_i uart.receive_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1678_ _0018_ clknet_4_8_0_wb_clk_i spi.div_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1063__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0980_ spi.div_counter\[3\] _0257_ spi.div_counter\[1\] spi.div_counter\[0\] _0379_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1532_ uart.div_counter\[4\] _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1601_ _0719_ _0815_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1394_ _0716_ _0699_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I RXD vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1463_ _0775_ _0778_ _0779_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1707__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0963_ _0284_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0894_ _0287_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1515_ _0819_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1377_ _0650_ _0706_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1446_ _0757_ _0762_ _0763_ _0764_ _0765_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1018__A1 spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1257__A1 _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1300_ uart.receive_div_counter\[4\] _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1162_ uart.receive_div_counter\[12\] uart.divisor\[12\] _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1231_ _0587_ _0588_ _0583_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1093_ _0468_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0877_ _0289_ _0291_ _0292_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0946_ spi.counter\[3\] _0339_ spi.counter\[4\] _0327_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1429_ _0749_ _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1411__A1 uart.div_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1780_ _0120_ clknet_4_5_0_wb_clk_i uart.div_counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1145_ _0459_ _0515_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1214_ _0567_ _0468_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1076_ net14 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0929_ _0330_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1632__A1 _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1694_ _0034_ clknet_4_12_0_wb_clk_i uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1763_ _0103_ clknet_4_1_0_wb_clk_i uart.data_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1059_ _0440_ _0434_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1128_ uart.divisor\[3\] _0462_ _0485_ spi.divisor\[3\] _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput25 net25 data_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1740__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0924__C _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1746_ _0086_ clknet_4_13_0_wb_clk_i uart.receive_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1677_ _0017_ clknet_4_8_0_wb_clk_i spi.div_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_15_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1763__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1462_ _0628_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1531_ _0816_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1600_ _0161_ _0204_ _0206_ _0248_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1393_ _0527_ _0538_ _0549_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1786__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1293__A2 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1729_ _0069_ clknet_4_3_0_wb_clk_i spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__0859__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0893_ _0271_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0962_ _0361_ _0364_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1514_ _0817_ _0815_ _0819_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1445_ _0247_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1376_ uart.receive_buff\[1\] _0702_ _0704_ uart.receive_buff\[2\] _0706_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_18_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1335__I _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1161_ uart.receive_div_counter\[9\] uart.divisor\[9\] _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1230_ uart.divisor\[13\] _0576_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1092_ _0425_ _0275_ _0463_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_47_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0945_ _0256_ _0270_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0876_ _0271_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1428_ uart.counter\[3\] uart.counter\[2\] _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1359_ _0690_ _0691_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_61_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1411__A2 uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1213_ _0432_ _0571_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1144_ _0497_ net23 _0514_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1075_ _0447_ _0452_ _0453_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0859_ _0275_ net2 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0928_ _0335_ _0334_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1396__A1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1594__B _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1148__B2 uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1693_ _0033_ clknet_4_12_0_wb_clk_i uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_40_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1762_ _0102_ clknet_4_0_0_wb_clk_i uart.data_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1127_ spi.dout\[3\] _0499_ _0469_ uart.divisor\[11\] _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1058_ net10 _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1692__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput26 net26 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_54_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0940__C _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1745_ _0085_ clknet_4_7_0_wb_clk_i uart.receive_div_counter\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ _0016_ clknet_4_8_0_wb_clk_i spi.div_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1392_ _0553_ _0700_ _0715_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1530_ _0144_ _0826_ _0147_ _0808_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1461_ _0776_ _0760_ _0777_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_45_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1728_ _0068_ clknet_4_3_0_wb_clk_i spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1730__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1659_ _0245_ _0246_ _0285_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_51_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0961_ _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1753__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0892_ _0297_ _0305_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1375_ _0650_ _0705_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1513_ uart.div_counter\[1\] _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1444_ _0754_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output26_I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1776__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1160_ uart.receive_div_counter\[14\] uart.divisor\[14\] _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1091_ _0425_ net3 _0463_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_55_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0944_ _0348_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_15_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0875_ net8 _0290_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1526__I uart.div_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1358_ uart.receive_div_counter\[13\] _0683_ _0682_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1427_ uart.counter\[1\] uart.counter\[0\] _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1799__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1289_ _0630_ _0631_ _0632_ _0633_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_38_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1166__A2 uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1212_ _0423_ _0571_ _0572_ _0574_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_47_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1143_ _0472_ _0511_ _0512_ _0513_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_35_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1074_ uart.divisor\[6\] _0445_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1081__I _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0927_ spi.counter\[0\] _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0858_ _0274_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1115__B _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1761_ _0101_ clknet_4_0_0_wb_clk_i uart.data_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1692_ _0032_ clknet_4_12_0_wb_clk_i uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1076__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1126_ _0474_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1057_ _0431_ _0438_ _0439_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput27 net27 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1302__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1744_ _0084_ clknet_4_5_0_wb_clk_i uart.receive_div_counter\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1675_ _0015_ clknet_4_10_0_wb_clk_i spi.div_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1109_ uart.divisor\[1\] _0462_ _0469_ uart.divisor\[9\] uart.dout\[1\] _0483_ _0484_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_51_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1039__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1391_ uart.receive_buff\[7\] _0704_ _0495_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1460_ _0773_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1303__B _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1682__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1658_ uart.dout\[7\] _0209_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1727_ _0067_ clknet_4_3_0_wb_clk_i spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1589_ _0191_ _0196_ _0197_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1439__I _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0960_ _0350_ _0328_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_54_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0891_ spi.data_out_buff\[2\] _0272_ _0304_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1512_ _0713_ _0818_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1374_ uart.receive_buff\[0\] _0702_ _0704_ uart.receive_buff\[1\] _0705_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1084__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1443_ _0757_ _0744_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1423__A1 uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1193__A3 _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1090_ uart.divisor\[0\] _0462_ _0465_ uart.dout\[0\] _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0943_ _0347_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1720__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0874_ _0278_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_15_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1288_ _0625_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1357_ uart.receive_div_counter\[14\] _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1426_ _0731_ _0743_ _0747_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1743__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1142_ uart.divisor\[5\] _0507_ _0479_ spi.divisor\[5\] _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1211_ _0573_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1073_ _0451_ _0433_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0857_ net3 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0926_ spi.counter\[1\] _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1409_ _0730_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_26_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1766__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1691_ _0031_ clknet_4_8_0_wb_clk_i net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1760_ _0100_ clknet_4_0_0_wb_clk_i uart.data_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1789__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1125_ uart.dout\[3\] _0483_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1056_ uart.divisor\[2\] _0428_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1267__I _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput28 net28 irq3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput17 net17 TXD vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_0909_ net13 _0314_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1743_ _0083_ clknet_4_7_0_wb_clk_i uart.receive_div_counter\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1087__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ _0014_ clknet_4_8_0_wb_clk_i spi.div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1108_ _0464_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1039_ net5 net6 _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1039__A2 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ _0713_ _0714_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1657_ uart.receive_buff\[7\] _0717_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1588_ _0191_ _0159_ _0194_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1726_ _0066_ clknet_4_2_0_wb_clk_i spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_48_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0890_ _0302_ _0303_ _0292_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1511_ _0812_ _0815_ _0817_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_10_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1442_ _0760_ _0761_ _0755_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1314__B _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1373_ _0703_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_61_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1709_ _0049_ clknet_4_15_0_wb_clk_i uart.receive_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1185__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1672__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0942_ net16 _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1405__A2 uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0873_ spi.data_out_buff\[1\] _0288_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1425_ _0744_ _0746_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1356_ _0687_ _0689_ _0673_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1341__A1 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1287_ _0630_ _0621_ uart.receive_div_counter\[0\] _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_50_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1695__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0902__I _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1141_ spi.dout\[5\] _0499_ _0505_ uart.divisor\[13\] _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1072_ net13 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1210_ _0283_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0856_ net4 _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_0925_ _0333_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1408_ _0720_ _0721_ _0724_ _0729_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_11_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1339_ uart.receive_div_counter\[10\] _0674_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1710__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1690_ _0030_ clknet_4_3_0_wb_clk_i spi.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1055_ _0437_ _0434_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1124_ _0460_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput18 net18 data_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_0839_ _0255_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0908_ spi.data_out_buff\[6\] _0307_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1283__I _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1742_ _0082_ clknet_4_5_0_wb_clk_i uart.receive_div_counter\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1673_ _0013_ clknet_4_8_0_wb_clk_i spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1756__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1107_ _0459_ _0482_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1038_ _0280_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1725_ _0065_ clknet_4_3_0_wb_clk_i spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1656_ _0243_ _0244_ _0285_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1587_ _0148_ _0195_ _0151_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_36_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1510_ _0812_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_10_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1441_ _0731_ _0743_ _0750_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1372_ _0552_ _0615_ _0616_ _0699_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1187__A2 _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1708_ _0048_ clknet_4_14_0_wb_clk_i net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1639_ _0230_ _0231_ _0232_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1178__A2 uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xserial_ports_30 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1102__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0941_ _0346_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_15_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0872_ _0287_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1355_ _0688_ _0683_ _0638_ _0682_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_50_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1424_ _0477_ _0745_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1286_ _0613_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1286__I _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1399__A2 uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1140_ uart.dout\[5\] _0465_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1071_ _0447_ _0449_ _0450_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_55_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0924_ _0249_ _0331_ _0292_ _0332_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_0855_ _0271_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1011__A1 spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1338_ _0638_ _0674_ uart.receive_div_counter\[10\] _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1407_ _0725_ _0726_ _0727_ _0728_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1269_ _0549_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1078__A1 uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1002__A1 _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1069__A1 _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1123_ _0491_ _0494_ _0496_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1054_ net9 _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1685__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1232__A1 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0907_ _0296_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput19 net19 data_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0838_ spi.divisor\[7\] _0250_ _0251_ spi.divisor\[4\] _0254_ _0255_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_19_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1741_ _0081_ clknet_4_7_0_wb_clk_i uart.receive_div_counter\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1672_ _0012_ clknet_4_8_0_wb_clk_i spi.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1106_ _0461_ net18 _0471_ _0481_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_48_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1037_ _0422_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1700__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1600__C _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1723__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1328__B _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1724_ _0064_ clknet_4_8_0_wb_clk_i spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1655_ uart.dout\[6\] _0237_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1586_ _0192_ _0194_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1746__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0831__I _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1371_ _0701_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_10_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1440_ _0759_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_61_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1707_ _0047_ clknet_4_15_0_wb_clk_i net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1638_ _0284_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1569_ _0180_ _0823_ _0173_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1769__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xserial_ports_31 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_55_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0940_ _0344_ _0331_ _0345_ _0337_ _0296_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__0861__A2 spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0871_ _0286_ spi.busy _0276_ _0277_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_2_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1354_ uart.receive_div_counter\[13\] _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1285_ uart.receive_div_counter\[2\] _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1423_ uart.busy _0277_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output17_I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1070_ uart.divisor\[5\] _0445_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0854_ _0249_ _0256_ _0270_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_0923_ _0247_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1337_ _0669_ _0664_ _0663_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1268_ _0538_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1406_ uart.div_counter\[7\] uart.divisor\[7\] _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1199_ _0550_ _0563_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_34_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1122_ _0461_ net20 _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1603__C _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1053_ _0431_ _0435_ _0436_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_38_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0837_ _0252_ spi.div_counter\[6\] spi.div_counter\[3\] _0253_ _0254_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_16_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0906_ _0297_ _0317_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input16_I rst vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1740_ _0080_ clknet_4_7_0_wb_clk_i uart.receive_div_counter\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1214__A2 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1671_ _0011_ clknet_4_10_0_wb_clk_i spi.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I data_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1105_ _0472_ _0480_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1036_ net26 _0396_ _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1141__B2 uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1675__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1435__A2 _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1199__A1 _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1654_ uart.receive_buff\[6\] _0235_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1723_ _0063_ clknet_4_9_0_wb_clk_i spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1585_ uart.div_counter\[8\] _0171_ _0193_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_0_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1019_ _0295_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1698__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1519__B _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1114__B2 spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1417__A2 uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1353__A1 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1370_ _0645_ _0700_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1637_ uart.dout\[1\] _0210_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1706_ _0046_ clknet_4_14_0_wb_clk_i net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1344__A1 _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1568_ _0178_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1499_ _0805_ _0798_ _0807_ _0808_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_36_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xserial_ports_32 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0870_ _0273_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1422_ uart.counter\[0\] _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1353_ _0631_ _0684_ uart.receive_div_counter\[13\] _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1284_ _0622_ _0627_ _0629_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1736__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0999_ _0335_ _0255_ _0269_ _0328_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_14_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0853_ _0269_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1759__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0922_ _0279_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_11_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1405_ uart.div_counter\[5\] uart.divisor\[5\] _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1336_ _0670_ _0672_ _0673_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1198_ uart.receive_counter\[1\] uart.receive_counter\[0\] uart.receive_counter\[2\]
+ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1267_ _0613_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput1 RXD net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1529__A1 uart.div_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1052_ uart.divisor\[1\] _0428_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1121_ _0347_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_31_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0836_ spi.divisor\[3\] _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0905_ spi.data_out_buff\[4\] _0306_ _0316_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1319_ uart.receive_div_counter\[7\] _0655_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1670_ _0010_ clknet_4_10_0_wb_clk_i spi.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1104_ spi.dout\[0\] _0475_ _0477_ uart.busy _0479_ spi.divisor\[0\] _0480_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_1035_ _0288_ _0363_ _0247_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1799_ _0139_ clknet_4_15_0_wb_clk_i uart.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_57_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_50_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ _0241_ _0242_ _0285_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1584_ uart.div_counter\[11\] uart.div_counter\[10\] uart.div_counter\[9\] _0193_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1722_ _0062_ clknet_4_9_0_wb_clk_i spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1018_ spi.dout\[3\] _0403_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1792__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0864__A1 _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1705_ _0045_ clknet_4_14_0_wb_clk_i net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1636_ uart.receive_buff\[1\] _0718_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1567_ _0178_ _0176_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1498_ _0573_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1665__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1023__A1 spi.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1421_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1352_ _0685_ _0686_ _0673_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1283_ _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1688__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1262__A1 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0998_ _0392_ _0393_ _0391_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1619_ spi.data_in_buff\[2\] _0218_ _0215_ spi.data_in_buff\[3\] _0220_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_37_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0921_ _0256_ _0270_ _0329_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_23_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0852_ _0259_ _0261_ _0265_ _0268_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1335_ _0628_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1404_ uart.div_counter\[4\] uart.divisor\[4\] _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1197_ _0561_ _0554_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1266_ uart.receiving _0553_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_36_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 addr[0] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1483__A1 _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1235__A1 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1226__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_27_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1009__I _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1051_ _0432_ _0434_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1120_ spi.divisor\[2\] _0485_ _0477_ uart.has_byte _0493_ _0494_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__1726__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0904_ _0313_ _0315_ _0310_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0835_ spi.divisor\[6\] _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1318_ _0656_ _0658_ _0629_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1249_ _0437_ _0599_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1749__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1150__A3 _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1103_ _0478_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1034_ _0418_ _0419_ _0420_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1610__A1 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1798_ _0138_ clknet_4_12_0_wb_clk_i uart.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1117__B1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1721_ _0061_ clknet_4_3_0_wb_clk_i uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_5_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1652_ uart.dout\[5\] _0237_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1583_ _0191_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1017_ spi.data_in_buff\[3\] _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1551__B _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0873__A2 _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0856__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1704_ _0044_ clknet_4_11_0_wb_clk_i net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1566_ uart.div_counter\[9\] _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1635_ _0228_ _0229_ _0190_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1497_ _0451_ _0794_ _0773_ _0806_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_36_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1351_ _0631_ _0684_ _0683_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1420_ _0736_ _0741_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1282_ _0283_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1210__I _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1366__B _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1618_ _0216_ _0219_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0997_ _0250_ _0376_ _0388_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_14_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1549_ _0159_ _0160_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1782__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0920_ _0328_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0851_ _0266_ _0267_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1334_ _0671_ _0626_ _0665_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1265_ uart.receive_div_counter\[0\] _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1403_ uart.div_counter\[13\] uart.divisor\[13\] _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1196_ uart.receive_counter\[3\] _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 addr[1] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_34_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0954__I _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_2_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1678__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1050_ _0433_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0834_ spi.div_counter\[4\] _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_0903_ net12 _0314_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1317_ _0651_ _0644_ _0657_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1248_ _0447_ _0600_ _0601_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1179_ uart.receive_div_counter\[3\] uart.divisor\[3\] _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1102_ _0286_ net3 _0463_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1033_ _0410_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1797_ _0137_ clknet_4_13_0_wb_clk_i uart.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input14_I data_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1117__A1 uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1117__B2 uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ uart.receive_buff\[5\] _0235_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1720_ _0060_ clknet_4_3_0_wb_clk_i uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1194__B _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1582_ uart.div_counter\[12\] _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I bus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1016_ _0329_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1739__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_31_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_61_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1634_ uart.dout\[0\] _0210_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1703_ _0043_ clknet_4_14_0_wb_clk_i net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1565_ _0175_ _0177_ _0169_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1496_ _0802_ _0799_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1350_ _0682_ _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1281_ _0623_ _0612_ _0626_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__0867__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0996_ spi.div_counter\[7\] _0389_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1617_ spi.data_in_buff\[1\] _0218_ _0215_ spi.data_in_buff\[2\] _0219_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1548_ uart.div_counter\[6\] _0162_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1479_ _0788_ _0781_ _0791_ _0792_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_37_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0850_ spi.divisor\[5\] spi.div_counter\[5\] _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1402_ _0722_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1333_ _0669_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1264_ _0610_ _0611_ _0593_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput4 addr[2] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1195_ _0558_ _0559_ _0560_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0979_ _0318_ _0378_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1171__A2 uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0880__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0833_ spi.div_counter\[7\] _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_0902_ _0278_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1772__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1316_ _0648_ _0654_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1178_ uart.receive_div_counter\[2\] uart.divisor\[2\] _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1247_ spi.divisor\[1\] _0595_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1126__I _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1795__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1101_ _0476_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1032_ spi.dout\[7\] _0402_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1796_ _0136_ clknet_4_12_0_wb_clk_i uart.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1668__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1650_ _0239_ _0240_ _0232_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_44_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1581_ _0188_ _0189_ _0190_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_53_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1015_ _0405_ _0406_ _0391_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1044__A1 uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1779_ _0119_ clknet_4_5_0_wb_clk_i uart.div_counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1035__A1 _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1274__A1 _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ uart.receive_buff\[0\] _0718_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1564_ uart.div_counter\[8\] _0176_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1702_ _0042_ clknet_4_14_0_wb_clk_i net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1495_ uart.data_buff\[8\] _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1280_ _0625_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1729__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0995_ _0387_ _0390_ _0391_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1547_ _0159_ _0160_ _0161_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1616_ _0395_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1478_ _0573_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1229__A1 _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1477__A1 _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1401_ uart.div_counter\[6\] uart.divisor\[6\] _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1194_ _0558_ _0559_ _0495_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1332_ _0669_ _0667_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1263_ spi.divisor\[7\] _0596_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput5 bus_cyc net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_34_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0978_ spi.div_counter\[3\] _0369_ _0376_ _0377_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1631__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0832_ spi.counter\[0\] _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0901_ spi.data_out_buff\[5\] _0307_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1315_ uart.receive_div_counter\[6\] _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1177_ uart.receive_div_counter\[4\] uart.divisor\[4\] _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1246_ _0432_ _0599_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1080__A2 _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1100_ net4 _0274_ _0473_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1031_ spi.data_in_buff\[7\] _0358_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1795_ _0135_ clknet_4_0_0_wb_clk_i net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_12_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1229_ _0448_ _0584_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1581__B _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1762__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1580_ _0284_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1014_ spi.dout\[2\] _0403_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1778_ _0118_ clknet_4_5_0_wb_clk_i uart.div_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1701_ _0041_ clknet_4_11_0_wb_clk_i net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1563_ _0148_ _0173_ _0161_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1632_ _0126_ _0227_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1494_ _0802_ _0798_ _0804_ _0792_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1505__I uart.div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0994_ _0356_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1546_ _0151_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1615_ _0216_ _0217_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1477_ _0437_ _0760_ _0789_ _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1410__A2 uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1401__A2 uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1331_ uart.receive_div_counter\[9\] _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1400_ uart.div_counter\[11\] uart.divisor\[11\] _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1193_ uart.receive_counter\[1\] uart.receive_counter\[0\] _0550_ _0559_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1262_ _0454_ _0603_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput6 bus_we net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_34_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0977_ _0262_ _0374_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1529_ uart.div_counter\[3\] _0814_ _0146_ _0827_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0900_ _0297_ _0312_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0831_ _0247_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1314_ _0618_ _0654_ _0645_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1176_ uart.receive_div_counter\[7\] uart.divisor\[7\] _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1245_ _0598_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1513__I uart.div_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_6_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1691__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0930__C _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1030_ _0416_ _0417_ _0411_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1794_ _0134_ clknet_4_2_0_wb_clk_i spi.data_in_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1228_ _0585_ _0586_ _0583_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1159_ uart.receiving _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1013_ spi.data_in_buff\[2\] _0359_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1777_ _0117_ clknet_4_5_0_wb_clk_i uart.div_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input12_I data_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1631_ net17 _0764_ _0226_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1700_ _0040_ clknet_4_10_0_wb_clk_i net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1562_ _0171_ _0174_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1493_ _0448_ _0794_ _0789_ _0803_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_1_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1752__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0993_ spi.div_counter\[6\] _0389_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1775__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1614_ spi.data_in_buff\[0\] _0396_ _0215_ spi.data_in_buff\[1\] _0217_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1183__A2 _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1545_ uart.div_counter\[6\] _0156_ _0150_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1476_ _0784_ _0785_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_59_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1174__A2 uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1798__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1330_ _0650_ _0668_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1165__A2 uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1261_ _0252_ _0595_ _0609_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1192_ uart.receive_counter\[2\] _0554_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 data_in[0] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0976_ _0363_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1528_ _0145_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1459_ uart.data_buff\[0\] _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0830_ net16 _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1313_ uart.receive_div_counter\[6\] _0651_ _0644_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_47_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1244_ _0567_ _0478_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_22_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1175_ _0539_ _0540_ _0541_ _0542_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__1074__A1 uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0959_ _0287_ _0329_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1065__A1 uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0879__A1 _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1056__A1 uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput10 data_in[3] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1793_ _0133_ clknet_4_0_0_wb_clk_i spi.data_in_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1709__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1158_ _0516_ _0526_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1227_ uart.divisor\[12\] _0577_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1089_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1012_ _0401_ _0404_ _0391_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1201__A1 _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _0116_ clknet_4_5_0_wb_clk_i uart.div_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1681__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0936__C _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1431__A1 _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1630_ _0776_ _0764_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1561_ _0154_ _0173_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1007__C _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1492_ _0797_ _0799_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1759_ _0099_ clknet_4_0_0_wb_clk_i uart.data_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1489__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0992_ _0350_ _0358_ _0388_ _0362_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1544_ _0816_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1613_ _0356_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1475_ _0772_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0921__A3 _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1191_ _0516_ _0557_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1260_ _0451_ _0596_ _0495_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput8 data_in[1] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1742__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0975_ _0263_ _0370_ _0375_ _0366_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1527_ uart.div_counter\[3\] _0825_ uart.div_counter\[1\] uart.div_counter\[0\] _0145_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1389_ uart.receive_buff\[6\] _0701_ _0709_ uart.receive_buff\[7\] _0714_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1458_ uart.data_buff\[1\] _0774_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1765__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1312_ _0650_ _0653_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_47_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1174_ uart.receive_div_counter\[5\] uart.divisor\[5\] _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1082__I _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1243_ _0423_ _0595_ _0597_ _0430_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0889_ net10 _0290_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0958_ spi.div_counter\[0\] _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1129__A3 _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0888__A2 _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1788__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 data_in[4] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1792_ _0132_ clknet_4_0_0_wb_clk_i spi.data_in_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1157_ net25 _0497_ _0525_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1226_ _0443_ _0584_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1088_ _0286_ _0275_ _0463_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_58_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1803__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1011_ spi.dout\[1\] _0403_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1775_ _0115_ clknet_4_5_0_wb_clk_i uart.div_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1209_ uart.divisor\[8\] _0570_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0951__A1 _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1445__I _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_53_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1560_ _0172_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1491_ uart.data_buff\[7\] _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1758_ _0098_ clknet_4_0_0_wb_clk_i uart.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1689_ _0029_ clknet_4_3_0_wb_clk_i spi.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xserial_ports_29 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_0_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1404__A2 uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0991_ _0260_ _0384_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_14_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1543_ _0713_ _0158_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1612_ _0213_ _0396_ _0215_ _0399_ _0765_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1671__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1474_ uart.data_buff\[4\] _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1034__B _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1694__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1190_ _0551_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_36_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 data_in[2] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0974_ _0257_ _0368_ _0363_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1526_ uart.div_counter\[3\] _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1457_ _0770_ _0768_ _0771_ _0774_ _0765_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_10_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1388_ _0356_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_56_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1311_ _0651_ _0646_ _0652_ _0626_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1543__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1173_ uart.receive_div_counter\[6\] uart.divisor\[6\] _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1242_ spi.divisor\[0\] _0596_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0888_ spi.data_out_buff\[3\] _0288_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0957_ _0357_ _0359_ _0360_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1206__C _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1534__A1 _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1509_ _0731_ _0743_ _0813_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_53_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1732__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1525__A1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0971__B _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput12 data_in[5] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1791_ _0131_ clknet_4_0_0_wb_clk_i spi.data_in_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1093__I _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1225_ _0570_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1156_ _0486_ _0522_ _0523_ _0524_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1087_ net2 _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1268__I _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1217__B _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1755__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1010_ _0402_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1778__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1774_ _0114_ clknet_4_4_0_wb_clk_i uart.div_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1208_ _0570_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1139_ _0459_ _0510_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1490_ _0797_ _0798_ _0801_ _0792_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_60_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1757_ _0097_ clknet_4_1_0_wb_clk_i uart.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1688_ _0028_ clknet_4_3_0_wb_clk_i spi.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I data_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1177__A2 uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0860__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1611_ _0214_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0990_ _0260_ _0382_ _0364_ _0383_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_14_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1168__A2 uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1542_ _0156_ _0152_ _0157_ _0823_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1473_ _0784_ _0781_ _0787_ _0574_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input2_I addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1398__A2 uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0842__A1 spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0973_ _0257_ _0367_ spi.div_counter\[0\] _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1387_ _0707_ _0712_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1525_ _0642_ _0828_ _0829_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_10_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1456_ _0773_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1077__A1 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1310_ _0651_ _0643_ _0640_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_47_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1241_ _0594_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1172_ uart.receive_div_counter\[8\] uart.divisor\[8\] _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1059__A1 _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0956_ spi.busy _0332_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0887_ _0297_ _0301_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1508_ _0814_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1439_ _0758_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1684__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput13 data_in[6] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_26_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1786__D _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1790_ _0130_ clknet_4_0_0_wb_clk_i spi.data_in_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1213__A1 _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1224_ _0581_ _0582_ _0583_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1086_ _0426_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1155_ uart.divisor\[7\] _0507_ _0479_ spi.divisor\[7\] _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0939_ _0344_ _0340_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1773_ _0113_ clknet_4_4_0_wb_clk_i uart.div_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1207_ _0424_ _0468_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1138_ _0497_ net22 _0509_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1069_ _0448_ _0433_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1722__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1745__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1099__I _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1756_ _0096_ clknet_4_0_0_wb_clk_i uart.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1687_ _0027_ clknet_4_2_0_wb_clk_i spi.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_13_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1768__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0860__A2 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1610_ _0278_ _0394_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1541_ _0156_ _0149_ _0146_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_1_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1472_ net8 _0760_ _0777_ _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_45_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1739_ _0079_ clknet_4_7_0_wb_clk_i uart.receive_div_counter\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1151__B _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0972_ _0371_ _0373_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1524_ _0819_ _0812_ _0825_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1386_ uart.receive_buff\[5\] _0701_ _0709_ uart.receive_buff\[6\] _0712_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1455_ _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1171_ uart.receive_div_counter\[0\] uart.divisor\[0\] _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1240_ _0594_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_56_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0886_ spi.data_out_buff\[1\] _0272_ _0300_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0955_ _0358_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1507_ _0759_ _0813_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1369_ _0615_ _0616_ _0699_ uart.receiving _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1438_ _0476_ _0745_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_53_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1289__A2 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput14 data_in[7] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1154_ spi.dout\[7\] _0475_ _0505_ uart.divisor\[15\] _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1223_ _0410_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1085_ _0460_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0869_ _0284_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0938_ spi.counter\[3\] _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1772_ _0112_ clknet_4_4_0_wb_clk_i uart.div_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1674__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1370__A1 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1137_ _0472_ _0504_ _0506_ _0508_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1206_ _0423_ _0568_ _0569_ _0366_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_18_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1068_ net12 _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1425__A2 _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1416__A2 uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1104__B2 uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1104__A1 spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1686_ _0026_ clknet_4_2_0_wb_clk_i spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1755_ _0095_ clknet_4_1_0_wb_clk_i uart.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1540_ uart.div_counter\[5\] _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_30_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0988__B _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1712__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1471_ _0780_ _0785_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1738_ _0078_ clknet_4_13_0_wb_clk_i uart.receive_div_counter\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1669_ _0009_ clknet_4_10_0_wb_clk_i spi.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1735__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0971_ _0367_ _0361_ _0372_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1523_ _0825_ _0815_ _0826_ _0827_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1454_ _0730_ _0742_ _0751_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1385_ _0707_ _0711_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1758__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output27_I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1170_ _0532_ _0537_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0885_ _0298_ _0299_ _0292_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0954_ _0329_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1437_ uart.counter\[1\] _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1506_ _0749_ _0750_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1368_ uart.receive_counter\[3\] _0563_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1299_ _0636_ _0632_ _0637_ _0641_ _0642_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_53_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 io_in net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1157__B _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1153_ uart.dout\[7\] _0465_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1222_ uart.divisor\[11\] _0577_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1084_ net5 _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0868_ _0283_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0937_ _0343_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1771_ _0111_ clknet_4_4_0_wb_clk_i uart.div_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1205_ uart_ien _0568_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1067_ _0348_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1136_ uart.divisor\[4\] _0507_ _0485_ spi.divisor\[4\] _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1260__B _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1754_ _0094_ clknet_4_13_0_wb_clk_i uart.receiving vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1791__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1685_ _0025_ clknet_4_2_0_wb_clk_i spi.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1119_ _0486_ _0492_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1664__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1470_ _0758_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1612__C _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1737_ _0077_ clknet_4_13_0_wb_clk_i uart.receive_div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1599_ _0827_ _0205_ uart.div_counter\[14\] _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1668_ _0008_ clknet_4_10_0_wb_clk_i spi.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1687__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1252__A1 _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0970_ _0347_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1243__A1 _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1522_ _0822_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1453_ uart.counter\[1\] _0744_ uart.counter\[2\] uart.counter\[3\] _0771_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1384_ uart.receive_buff\[4\] _0701_ _0709_ uart.receive_buff\[5\] _0711_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1216__A1 uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0884_ net9 _0290_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0953_ _0356_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1367_ _0696_ _0697_ _0698_ _0574_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1505_ uart.div_counter\[0\] _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1436_ _0756_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1298_ _0573_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1725__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1207__A1 _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput16 rst net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1221_ _0440_ _0571_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_9_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1748__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1152_ _0516_ _0521_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1083_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0936_ _0339_ _0331_ _0342_ _0337_ _0332_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_7_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0867_ net16 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1419_ _0737_ _0738_ _0739_ _0740_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1770_ _0110_ clknet_4_4_0_wb_clk_i uart.div_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1204_ _0567_ _0467_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1066_ _0431_ _0444_ _0446_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1135_ _0426_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0919_ spi.counter\[3\] spi.counter\[2\] spi.counter\[4\] _0327_ _0328_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_7_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1451__B _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1753_ _0093_ clknet_4_13_0_wb_clk_i uart.receive_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ _0024_ clknet_4_2_0_wb_clk_i spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1118_ spi.dout\[2\] _0475_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1049_ _0425_ _0276_ _0277_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_50_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1736_ _0076_ clknet_4_13_0_wb_clk_i uart.receive_div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_17_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1598_ _0194_ _0203_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1667_ _0007_ clknet_4_10_0_wb_clk_i spi.data_out_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1781__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1383_ _0707_ _0710_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1521_ _0825_ _0819_ uart.div_counter\[0\] _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1452_ uart.counter\[3\] _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1719_ _0059_ clknet_4_6_0_wb_clk_i uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0952_ _0283_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0883_ spi.data_out_buff\[2\] _0288_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1677__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1504_ _0809_ _0768_ _0774_ _0808_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1152__A1 _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1366_ _0633_ _0693_ _0613_ _0696_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_10_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1435_ _0748_ _0126_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1297_ _0638_ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_43_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1207__A2 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_61_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1151_ _0461_ net24 _0520_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1220_ _0579_ _0580_ _0420_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1134__A1 spi.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1082_ _0295_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0866_ _0248_ _0272_ _0282_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_23_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0935_ _0340_ _0341_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1349_ _0683_ _0682_ _0617_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1418_ uart.div_counter\[0\] uart.divisor\[0\] _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1539__B _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1715__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1134_ spi.dout\[4\] _0499_ _0505_ uart.divisor\[12\] _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1203_ _0424_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1065_ uart.divisor\[4\] _0445_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1203__I _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0918_ spi.counter\[0\] spi.counter\[1\] _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0849_ spi.divisor\[1\] spi.div_counter\[1\] _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0952__I _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1738__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_60_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0862__I _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1752_ _0092_ clknet_4_15_0_wb_clk_i uart.receive_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _0023_ clknet_4_8_0_wb_clk_i spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1117_ uart.divisor\[2\] _0462_ _0469_ uart.divisor\[10\] uart.dout\[2\] _0483_ _0491_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_0_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1048_ net8 _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_8_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1446__C _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0857__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1735_ _0075_ clknet_4_13_0_wb_clk_i uart.receive_div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1666_ _0006_ clknet_4_10_0_wb_clk_i spi.data_out_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1597_ _0202_ _0194_ _0203_ _0822_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1520_ uart.div_counter\[2\] _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1382_ uart.receive_buff\[3\] _0702_ _0709_ uart.receive_buff\[4\] _0710_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1451_ _0767_ _0769_ _0642_ _0752_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_26_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1649_ uart.dout\[4\] _0237_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1718_ _0058_ clknet_4_6_0_wb_clk_i uart.divisor\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1161__A2 uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_55_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0882_ _0296_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0951_ _0349_ _0353_ _0354_ _0355_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_12_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1503_ _0809_ _0798_ _0811_ _0808_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1296_ _0639_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1365_ _0690_ _0633_ _0691_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1434_ _0744_ _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0966__A2 _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1771__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1150_ _0486_ _0517_ _0518_ _0519_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_9_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1081_ _0457_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1070__A1 uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0865_ spi.data_out_buff\[0\] _0279_ _0281_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_21_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1794__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0934_ _0249_ _0334_ _0339_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1417_ uart.div_counter\[8\] uart.divisor\[8\] _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1279_ _0552_ _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1348_ uart.receive_div_counter\[12\] _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1667__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0875__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1052__A1 uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1202_ _0566_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1064_ _0427_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1133_ _0468_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__0866__A1 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1291__A1 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0917_ _0318_ _0326_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0848_ spi.divisor\[3\] _0262_ _0263_ spi.divisor\[2\] _0264_ _0265_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0848__A1 spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _0091_ clknet_4_15_0_wb_clk_i uart.receive_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1682_ _0022_ clknet_4_8_0_wb_clk_i net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1116_ _0484_ _0489_ _0490_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1047_ _0348_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1255__A1 spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1803_ _0143_ clknet_4_15_0_wb_clk_i uart.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1246__A1 _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1734_ _0074_ clknet_4_7_0_wb_clk_i uart.receive_div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1596_ uart.div_counter\[13\] _0191_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ _0005_ clknet_4_10_0_wb_clk_i spi.data_out_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1653__B _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1728__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1457__C _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1450_ _0731_ _0743_ _0768_ uart.counter\[2\] _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1381_ _0703_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0868__I _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1219__A1 uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1367__C _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1648_ uart.receive_buff\[4\] _0235_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1579_ uart.div_counter\[11\] _0183_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1717_ _0057_ clknet_4_6_0_wb_clk_i uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0881_ _0295_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0950_ _0256_ _0270_ _0279_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1433_ _0730_ _0742_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1502_ _0454_ _0785_ _0773_ _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1295_ uart.receive_div_counter\[3\] _0630_ uart.receive_div_counter\[1\] uart.receive_div_counter\[0\]
+ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1364_ uart.receive_div_counter\[15\] _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1612__A1 _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1143__A3 _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1080_ uart_ien _0349_ uart.has_byte _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0881__I _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0864_ _0280_ _0279_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0933_ _0249_ _0334_ _0339_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1347_ _0643_ _0639_ _0662_ _0681_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1416_ uart.div_counter\[10\] uart.divisor\[10\] _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1278_ _0615_ _0616_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1201_ _0349_ _0565_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1132_ uart.dout\[4\] _0483_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1063_ _0443_ _0434_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1761__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0916_ spi.data_out_buff\[6\] _0306_ _0325_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1656__B _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0847_ spi.divisor\[0\] spi.div_counter\[0\] _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1391__B _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1784__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ _0090_ clknet_4_15_0_wb_clk_i uart.receive_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _0021_ clknet_4_2_0_wb_clk_i spi.div_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I data_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1115_ _0461_ net19 _0372_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1046_ _0423_ _0428_ _0429_ _0430_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_39_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1191__A1 _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1733_ _0073_ clknet_4_6_0_wb_clk_i uart.receive_div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1802_ _0142_ clknet_4_14_0_wb_clk_i uart.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1595_ uart.div_counter\[14\] _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1664_ _0004_ clknet_4_10_0_wb_clk_i spi.data_out_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1029_ spi.dout\[6\] _0402_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1380_ _0707_ _0708_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1473__C _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1716_ _0056_ clknet_4_6_0_wb_clk_i uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_5_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1647_ _0236_ _0238_ _0232_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1578_ _0182_ _0187_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1155__A1 uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1155__B2 spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0880_ net16 _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_30_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1468__C _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1363_ _0694_ _0695_ _0673_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1432_ _0753_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1501_ _0805_ _0799_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1294_ _0625_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1659__B _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1128__A1 uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1128__B2 spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0932_ spi.counter\[2\] _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0863_ net7 _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__1690__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1346_ uart.receive_div_counter\[11\] uart.receive_div_counter\[10\] _0669_ _0664_
+ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1415_ uart.div_counter\[14\] uart.divisor\[14\] _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1277_ _0621_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1200_ _0562_ _0564_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1512__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1131_ _0459_ _0503_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1062_ net11 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1002__B net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0915_ _0323_ _0324_ _0310_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0846_ spi.div_counter\[2\] _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1329_ _0663_ _0666_ _0667_ _0664_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1048__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ _0020_ clknet_4_2_0_wb_clk_i spi.div_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1114_ spi.divisor\[1\] _0485_ _0477_ spi.busy _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1045_ _0348_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1421__I _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1751__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1732_ _0072_ clknet_4_13_0_wb_clk_i uart.receive_div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1801_ _0141_ clknet_4_14_0_wb_clk_i uart.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1663_ _0003_ clknet_4_11_0_wb_clk_i spi.data_out_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1182__A2 _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1594_ _0199_ _0201_ _0190_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1028_ spi.data_in_buff\[6\] _0407_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1774__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1173__A2 uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1646_ uart.dout\[3\] _0237_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1715_ _0055_ clknet_4_12_0_wb_clk_i uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1577_ uart.div_counter\[11\] _0154_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1146__I _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1500_ uart.data_buff\[9\] _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1362_ _0690_ _0614_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1293_ uart.receive_div_counter\[3\] _0631_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1431_ _0295_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1073__A1 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1629_ _0357_ _0225_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1055__A1 _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0931_ _0338_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0862_ _0278_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1276_ _0619_ _0614_ _0621_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1345_ uart.receive_div_counter\[11\] _0677_ _0680_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1414_ _0732_ _0733_ _0734_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1046__A1 _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1299__C _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1130_ _0497_ net21 _0502_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_25_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1061_ _0431_ _0441_ _0442_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_34_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0845_ spi.div_counter\[3\] _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_0914_ net14 _0314_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1328_ _0618_ _0665_ _0645_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1259_ _0607_ _0608_ _0593_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1680__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1044_ uart.divisor\[0\] _0427_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1113_ _0486_ _0487_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1497__A1 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1249__A1 _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_39_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1412__A1 uart.div_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1800_ _0140_ clknet_4_14_0_wb_clk_i uart.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ _0071_ clknet_4_7_0_wb_clk_i uart.receive_div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1662_ _0002_ clknet_4_11_0_wb_clk_i spi.data_out_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1593_ _0195_ _0200_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_28_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1027_ _0414_ _0415_ _0411_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_42_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1645_ _0209_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1576_ _0184_ _0186_ _0169_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1714_ _0054_ clknet_4_12_0_wb_clk_i uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1741__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1091__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1606__A1 _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1430_ _0751_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1361_ _0638_ _0692_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1292_ uart.receive_div_counter\[3\] _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1137__A3 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1764__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1559_ uart.div_counter\[8\] _0171_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1628_ spi.data_in_buff\[6\] _0395_ _0221_ spi.data_in_buff\[7\] _0225_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1787__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0861_ _0273_ spi.busy _0276_ _0277_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_0930_ _0334_ _0331_ _0336_ _0337_ _0332_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1413_ uart.div_counter\[12\] uart.divisor\[12\] _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1344_ _0372_ _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1275_ uart.receive_div_counter\[1\] _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1521__A3 uart.div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_0_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1060_ uart.divisor\[3\] _0428_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0913_ spi.data_out_buff\[7\] _0307_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0844_ spi.divisor\[6\] _0260_ _0251_ spi.divisor\[4\] _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1327_ _0648_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1189_ uart.receive_counter\[1\] _0554_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1258_ spi.divisor\[5\] _0596_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1043_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1112_ spi.dout\[1\] _0475_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input15_I io_in vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1412__A2 uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1100__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1730_ _0070_ clknet_4_13_0_wb_clk_i uart.receive_div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_40_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1592_ uart.div_counter\[13\] _0154_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1403__A2 uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1661_ _0001_ clknet_4_11_0_wb_clk_i spi.data_out_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input7_I data_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0914__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1026_ spi.dout\[5\] _0402_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1158__A1 _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1670__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1094__B1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1149__A1 uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1713_ _0053_ clknet_4_11_0_wb_clk_i uart_ien vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1644_ uart.receive_buff\[3\] _0235_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1575_ _0178_ _0173_ _0185_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1693__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1009_ _0351_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1360_ _0690_ _0691_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1291_ _0248_ _0634_ _0635_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1558_ _0149_ _0145_ _0170_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1627_ _0357_ _0224_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1489_ _0443_ _0794_ _0789_ _0800_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_17_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1122__B _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0860_ net5 net6 _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_2_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1343_ _0648_ _0676_ _0678_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1731__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1083__I _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1412_ uart.div_counter\[3\] uart.divisor\[3\] _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1274_ _0516_ _0620_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0989_ _0385_ _0386_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_57_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1754__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0912_ _0318_ _0322_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1036__I0 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0843_ spi.div_counter\[6\] _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1326_ _0664_ _0663_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1188_ _0551_ _0555_ _0420_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1257_ _0448_ _0603_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1777__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1042_ _0424_ _0426_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1111_ _0460_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1309_ uart.receive_div_counter\[5\] _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1271__I _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1220__B _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1176__A2 uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1591_ uart.div_counter\[13\] _0196_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1660_ _0000_ clknet_4_11_0_wb_clk_i spi.data_out_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_46_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1025_ spi.data_in_buff\[5\] _0407_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_55_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1789_ _0129_ clknet_4_2_0_wb_clk_i spi.data_in_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1094__B2 uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1712_ _0052_ clknet_4_15_0_wb_clk_i uart.receive_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1643_ _0717_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1574_ _0159_ _0182_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1035__B _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1008_ spi.data_in_buff\[1\] _0359_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1290_ _0621_ _0612_ _0630_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_46_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1230__A1 uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1626_ spi.data_in_buff\[5\] _0395_ _0221_ spi.data_in_buff\[6\] _0224_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1557_ uart.div_counter\[7\] uart.div_counter\[6\] uart.div_counter\[5\] _0170_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1488_ _0793_ _0799_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1212__C _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1221__A1 _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1683__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1212__A1 _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1342_ uart.receive_div_counter\[11\] _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1273_ _0612_ _0614_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1411_ uart.div_counter\[1\] uart.divisor\[1\] _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0988_ _0382_ _0383_ _0372_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1609_ net15 _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1449__I _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0911_ spi.data_out_buff\[5\] _0306_ _0321_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0842_ spi.divisor\[7\] _0250_ _0257_ _0258_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_59_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1325_ uart.receive_div_counter\[8\] _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1256_ _0605_ _0606_ _0593_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1187_ uart.receive_counter\[0\] _0550_ _0554_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1721__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1110_ _0478_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1041_ _0425_ _0276_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1308_ _0458_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1744__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1239_ _0567_ _0478_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1462__I _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1590_ _0713_ _0198_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1024_ _0412_ _0413_ _0411_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1767__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1788_ _0128_ clknet_4_2_0_wb_clk_i spi.data_in_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1282__I _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0964__C _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1711_ _0051_ clknet_4_15_0_wb_clk_i uart.receive_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1642_ _0233_ _0234_ _0232_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1573_ uart.div_counter\[10\] _0183_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1007_ _0399_ _0359_ _0400_ _0366_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_16_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_32_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1097__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1556_ _0166_ _0168_ _0169_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1625_ _0357_ _0223_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1487_ _0759_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_32_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1470__I _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1410_ uart.div_counter\[9\] uart.divisor\[9\] _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1272_ _0612_ _0618_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1341_ _0248_ _0675_ _0677_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_46_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0987_ _0382_ _0369_ _0364_ _0384_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1555__I _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1608_ _0210_ _0212_ _0190_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1539_ _0153_ _0155_ _0779_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_57_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_19_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0910_ _0319_ _0320_ _0310_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0841_ spi.divisor\[2\] _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1433__A2 _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1324_ _0643_ _0639_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1186_ _0552_ _0553_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1255_ spi.divisor\[4\] _0595_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1673__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1112__A1 spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1415__A2 uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1351__A1 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1040_ net4 _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1406__A2 uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1696__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1590__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1307_ _0647_ _0649_ _0629_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1169_ _0533_ _0534_ _0535_ _0536_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_1238_ _0591_ _0592_ _0593_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1023_ spi.dout\[4\] _0403_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1787_ _0127_ clknet_4_2_0_wb_clk_i spi.data_in_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1711__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input13_I data_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0907__I _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1734__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1710_ _0050_ clknet_4_15_0_wb_clk_i uart.receive_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1641_ uart.dout\[2\] _0210_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1572_ _0148_ _0182_ _0161_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I bus_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1006_ spi.dout\[0\] _0358_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1527__A1 uart.div_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1757__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0975__C _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1378__I _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1555_ _0628_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1624_ spi.data_in_buff\[4\] _0218_ _0221_ spi.data_in_buff\[5\] _0223_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1486_ _0777_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1340_ _0633_ _0676_ _0613_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0830__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1271_ _0617_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0986_ _0382_ _0383_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1607_ uart.has_byte _0211_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1538_ uart.div_counter\[4\] _0154_ _0146_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1469_ uart.data_buff\[3\] _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0840_ spi.div_counter\[2\] _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1323_ uart.receive_div_counter\[7\] uart.receive_div_counter\[6\] uart.receive_div_counter\[5\]
+ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_51_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1185_ net1 _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1254_ _0443_ _0603_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_20_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1340__B _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0969_ _0367_ _0369_ _0364_ _0370_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1179__A2 uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1306_ uart.receive_div_counter\[4\] _0648_ _0640_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1168_ uart.receive_div_counter\[15\] uart.divisor\[15\] _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1099_ _0474_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1237_ _0410_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1790__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0844__B2 spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1022_ spi.data_in_buff\[4\] _0407_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1260__A1 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1786_ _0126_ clknet_4_1_0_wb_clk_i uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0923__I _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_42_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1686__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1640_ uart.receive_buff\[2\] _0718_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1571_ uart.div_counter\[10\] _0178_ _0172_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_49_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1005_ spi.data_in_buff\[0\] _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1233__A1 uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1769_ _0109_ clknet_4_4_0_wb_clk_i uart.div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1472__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1608__B _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1554_ _0167_ _0823_ _0160_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1623_ _0216_ _0222_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1485_ uart.data_buff\[6\] _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
.ends

